
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity OSDBoot_ROM is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of OSDBoot_ROM is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"01",x"c9",x"87",x"04"),
     1 => (x"cc",x"87",x"03",x"cf"),
     2 => (x"87",x"00",x"fd",x"87"),
     3 => (x"27",x"29",x"00",x"00"),
     4 => (x"00",x"4f",x"27",x"36"),
     5 => (x"00",x"00",x"00",x"4f"),
     6 => (x"0e",x"18",x"1e",x"0e"),
     7 => (x"27",x"44",x"00",x"00"),
     8 => (x"00",x"0f",x"26",x"48"),
     9 => (x"ff",x"80",x"26",x"08"),
    10 => (x"4f",x"c0",x"e0",x"c0"),
    11 => (x"4e",x"27",x"f9",x"02"),
    12 => (x"00",x"00",x"0f",x"00"),
    13 => (x"fd",x"87",x"c0",x"d0"),
    14 => (x"c0",x"4e",x"27",x"43"),
    15 => (x"00",x"00",x"00",x"0f"),
    16 => (x"00",x"fd",x"87",x"4f"),
    17 => (x"0e",x"18",x"1e",x"0e"),
    18 => (x"26",x"48",x"ff",x"80"),
    19 => (x"26",x"08",x"4f",x"0e"),
    20 => (x"5e",x"5a",x"5b",x"5c"),
    21 => (x"5d",x"0e",x"1e",x"d8"),
    22 => (x"66",x"4d",x"76",x"49"),
    23 => (x"c0",x"79",x"75",x"49"),
    24 => (x"c0",x"b7",x"a9",x"03"),
    25 => (x"c0",x"ce",x"87",x"c0"),
    26 => (x"ed",x"1e",x"27",x"a6"),
    27 => (x"14",x"00",x"00",x"0f"),
    28 => (x"c4",x"86",x"c0",x"0d"),
    29 => (x"8d",x"75",x"9d",x"02"),
    30 => (x"c1",x"c6",x"87",x"c0"),
    31 => (x"4c",x"75",x"4a",x"dc"),
    32 => (x"b7",x"2a",x"72",x"4b"),
    33 => (x"cf",x"9b",x"c4",x"35"),
    34 => (x"73",x"9b",x"02",x"c0"),
    35 => (x"c4",x"87",x"76",x"49"),
    36 => (x"c1",x"79",x"73",x"49"),
    37 => (x"c9",x"b7",x"a9",x"06"),
    38 => (x"c0",x"c6",x"87",x"c0"),
    39 => (x"f7",x"83",x"c0",x"c3"),
    40 => (x"87",x"c0",x"f0",x"83"),
    41 => (x"6e",x"02",x"c0",x"ca"),
    42 => (x"87",x"73",x"1e",x"27"),
    43 => (x"a6",x"14",x"00",x"00"),
    44 => (x"0f",x"c4",x"86",x"c1"),
    45 => (x"84",x"74",x"49",x"c8"),
    46 => (x"b7",x"a9",x"04",x"fe"),
    47 => (x"ff",x"87",x"c0",x"cb"),
    48 => (x"87",x"c0",x"f0",x"1e"),
    49 => (x"27",x"a6",x"14",x"00"),
    50 => (x"00",x"0f",x"c4",x"86"),
    51 => (x"c0",x"48",x"26",x"26"),
    52 => (x"4d",x"26",x"4c",x"26"),
    53 => (x"4b",x"26",x"4a",x"26"),
    54 => (x"4f",x"0e",x"5e",x"5a"),
    55 => (x"5b",x"5c",x"5d",x"0e"),
    56 => (x"1e",x"c0",x"4c",x"76"),
    57 => (x"49",x"c0",x"79",x"dc"),
    58 => (x"a6",x"4b",x"d8",x"66"),
    59 => (x"4a",x"d8",x"66",x"48"),
    60 => (x"c1",x"80",x"dc",x"a6"),
    61 => (x"58",x"12",x"4d",x"d8"),
    62 => (x"35",x"b7",x"2d",x"75"),
    63 => (x"9d",x"02",x"c4",x"d7"),
    64 => (x"87",x"6e",x"02",x"c3"),
    65 => (x"e1",x"87",x"76",x"49"),
    66 => (x"c0",x"79",x"75",x"4a"),
    67 => (x"75",x"49",x"c1",x"e3"),
    68 => (x"a9",x"02",x"c2",x"e5"),
    69 => (x"87",x"72",x"49",x"c1"),
    70 => (x"e4",x"a9",x"02",x"c0"),
    71 => (x"de",x"87",x"72",x"49"),
    72 => (x"c1",x"ec",x"a9",x"02"),
    73 => (x"c2",x"cc",x"87",x"72"),
    74 => (x"49",x"c1",x"f3",x"a9"),
    75 => (x"02",x"c1",x"ea",x"87"),
    76 => (x"72",x"49",x"c1",x"f8"),
    77 => (x"a9",x"02",x"c0",x"f2"),
    78 => (x"87",x"c2",x"d3",x"87"),
    79 => (x"ca",x"1e",x"27",x"40"),
    80 => (x"18",x"00",x"00",x"1e"),
    81 => (x"c4",x"83",x"73",x"4a"),
    82 => (x"c4",x"8a",x"6a",x"1e"),
    83 => (x"27",x"4f",x"00",x"00"),
    84 => (x"00",x"0f",x"cc",x"86"),
    85 => (x"70",x"4a",x"74",x"4c"),
    86 => (x"72",x"84",x"27",x"40"),
    87 => (x"18",x"00",x"00",x"1e"),
    88 => (x"27",x"b5",x"14",x"00"),
    89 => (x"00",x"0f",x"c4",x"86"),
    90 => (x"c2",x"d6",x"87",x"d0"),
    91 => (x"1e",x"27",x"40",x"18"),
    92 => (x"00",x"00",x"1e",x"c4"),
    93 => (x"83",x"73",x"4a",x"c4"),
    94 => (x"8a",x"6a",x"1e",x"27"),
    95 => (x"4f",x"00",x"00",x"00"),
    96 => (x"0f",x"cc",x"86",x"70"),
    97 => (x"4a",x"74",x"4c",x"72"),
    98 => (x"84",x"27",x"40",x"18"),
    99 => (x"00",x"00",x"1e",x"27"),
   100 => (x"b5",x"14",x"00",x"00"),
   101 => (x"0f",x"c4",x"86",x"c1"),
   102 => (x"e7",x"87",x"c4",x"83"),
   103 => (x"73",x"4a",x"c4",x"8a"),
   104 => (x"6a",x"1e",x"27",x"b5"),
   105 => (x"14",x"00",x"00",x"0f"),
   106 => (x"c4",x"86",x"70",x"4a"),
   107 => (x"74",x"4c",x"72",x"84"),
   108 => (x"c1",x"ce",x"87",x"76"),
   109 => (x"49",x"c1",x"79",x"c1"),
   110 => (x"c7",x"87",x"c4",x"83"),
   111 => (x"73",x"4a",x"c4",x"8a"),
   112 => (x"6a",x"1e",x"27",x"a6"),
   113 => (x"14",x"00",x"00",x"0f"),
   114 => (x"c4",x"86",x"c1",x"84"),
   115 => (x"c0",x"f2",x"87",x"c0"),
   116 => (x"e5",x"1e",x"27",x"a6"),
   117 => (x"14",x"00",x"00",x"0f"),
   118 => (x"c4",x"86",x"75",x"1e"),
   119 => (x"27",x"a6",x"14",x"00"),
   120 => (x"00",x"0f",x"c4",x"86"),
   121 => (x"c0",x"da",x"87",x"75"),
   122 => (x"49",x"c0",x"e5",x"a9"),
   123 => (x"05",x"c0",x"c7",x"87"),
   124 => (x"76",x"49",x"c1",x"79"),
   125 => (x"c0",x"ca",x"87",x"75"),
   126 => (x"1e",x"27",x"a6",x"14"),
   127 => (x"00",x"00",x"0f",x"c4"),
   128 => (x"86",x"d8",x"66",x"4a"),
   129 => (x"d8",x"66",x"48",x"c1"),
   130 => (x"80",x"dc",x"a6",x"58"),
   131 => (x"12",x"4d",x"d8",x"35"),
   132 => (x"b7",x"2d",x"75",x"9d"),
   133 => (x"05",x"fb",x"e9",x"87"),
   134 => (x"74",x"48",x"26",x"26"),
   135 => (x"4d",x"26",x"4c",x"26"),
   136 => (x"4b",x"26",x"4a",x"26"),
   137 => (x"4f",x"0e",x"5e",x"5a"),
   138 => (x"5b",x"0e",x"cc",x"66"),
   139 => (x"4a",x"d8",x"b7",x"2a"),
   140 => (x"c3",x"ff",x"9a",x"cc"),
   141 => (x"66",x"4b",x"c8",x"b7"),
   142 => (x"2b",x"cf",x"fc",x"c0"),
   143 => (x"9b",x"72",x"4a",x"73"),
   144 => (x"b2",x"cc",x"66",x"4b"),
   145 => (x"c8",x"33",x"c0",x"ff"),
   146 => (x"f0",x"c0",x"c0",x"9b"),
   147 => (x"72",x"4a",x"73",x"b2"),
   148 => (x"cc",x"66",x"4b",x"d8"),
   149 => (x"33",x"cf",x"fc",x"c0"),
   150 => (x"c0",x"c0",x"9b",x"72"),
   151 => (x"4a",x"73",x"b2",x"72"),
   152 => (x"48",x"26",x"4b",x"26"),
   153 => (x"4a",x"26",x"4f",x"0e"),
   154 => (x"5e",x"5a",x"5b",x"0e"),
   155 => (x"cc",x"66",x"4a",x"c8"),
   156 => (x"b7",x"2a",x"c3",x"ff"),
   157 => (x"9a",x"cc",x"66",x"4b"),
   158 => (x"c8",x"33",x"cf",x"fc"),
   159 => (x"c0",x"9b",x"72",x"4a"),
   160 => (x"73",x"b2",x"72",x"48"),
   161 => (x"26",x"4b",x"26",x"4a"),
   162 => (x"26",x"4f",x"0e",x"5e"),
   163 => (x"5a",x"5b",x"0e",x"cc"),
   164 => (x"66",x"4a",x"d0",x"b7"),
   165 => (x"2a",x"cf",x"ff",x"ff"),
   166 => (x"9a",x"4a",x"cc",x"66"),
   167 => (x"4b",x"d0",x"33",x"f0"),
   168 => (x"c0",x"c0",x"9b",x"72"),
   169 => (x"4a",x"73",x"b2",x"72"),
   170 => (x"48",x"26",x"4b",x"26"),
   171 => (x"4a",x"26",x"4f",x"0e"),
   172 => (x"5e",x"5a",x"5b",x"5c"),
   173 => (x"5d",x"0e",x"d8",x"66"),
   174 => (x"4d",x"c0",x"4c",x"d4"),
   175 => (x"66",x"4a",x"dc",x"b7"),
   176 => (x"2a",x"72",x"4b",x"cf"),
   177 => (x"9b",x"d4",x"66",x"48"),
   178 => (x"c4",x"30",x"d8",x"a6"),
   179 => (x"58",x"73",x"49",x"c9"),
   180 => (x"b7",x"a9",x"06",x"c0"),
   181 => (x"c6",x"87",x"c0",x"f7"),
   182 => (x"83",x"c0",x"c3",x"87"),
   183 => (x"c0",x"f0",x"83",x"73"),
   184 => (x"97",x"7d",x"c1",x"85"),
   185 => (x"c1",x"84",x"74",x"49"),
   186 => (x"c8",x"b7",x"a9",x"04"),
   187 => (x"ff",x"cc",x"87",x"26"),
   188 => (x"4d",x"26",x"4c",x"26"),
   189 => (x"4b",x"26",x"4a",x"26"),
   190 => (x"4f",x"0e",x"5e",x"5a"),
   191 => (x"5b",x"5c",x"5d",x"0e"),
   192 => (x"cc",x"8e",x"27",x"26"),
   193 => (x"16",x"00",x"00",x"1e"),
   194 => (x"27",x"9e",x"0d",x"00"),
   195 => (x"00",x"0f",x"c4",x"86"),
   196 => (x"27",x"3c",x"16",x"00"),
   197 => (x"00",x"1e",x"27",x"b5"),
   198 => (x"14",x"00",x"00",x"0f"),
   199 => (x"c4",x"86",x"27",x"f5"),
   200 => (x"12",x"00",x"00",x"0f"),
   201 => (x"c0",x"86",x"70",x"4a"),
   202 => (x"72",x"9a",x"02",x"c4"),
   203 => (x"fd",x"87",x"27",x"0f"),
   204 => (x"16",x"00",x"00",x"1e"),
   205 => (x"27",x"b5",x"14",x"00"),
   206 => (x"00",x"0f",x"c4",x"86"),
   207 => (x"27",x"dc",x"04",x"00"),
   208 => (x"00",x"0f",x"c0",x"86"),
   209 => (x"70",x"4a",x"72",x"9a"),
   210 => (x"02",x"c4",x"c0",x"87"),
   211 => (x"27",x"00",x"20",x"00"),
   212 => (x"00",x"bf",x"1e",x"27"),
   213 => (x"b6",x"15",x"00",x"00"),
   214 => (x"1e",x"27",x"0b",x"0c"),
   215 => (x"00",x"00",x"0f",x"c8"),
   216 => (x"86",x"70",x"4b",x"73"),
   217 => (x"9b",x"02",x"c3",x"d2"),
   218 => (x"87",x"c4",x"a6",x"49"),
   219 => (x"27",x"00",x"20",x"00"),
   220 => (x"00",x"79",x"c0",x"4d"),
   221 => (x"c3",x"83",x"fc",x"9b"),
   222 => (x"27",x"00",x"20",x"00"),
   223 => (x"00",x"bf",x"4c",x"73"),
   224 => (x"84",x"74",x"1e",x"27"),
   225 => (x"aa",x"15",x"00",x"00"),
   226 => (x"1e",x"27",x"0b",x"0c"),
   227 => (x"00",x"00",x"0f",x"c8"),
   228 => (x"86",x"70",x"4a",x"72"),
   229 => (x"9a",x"02",x"c3",x"e0"),
   230 => (x"87",x"73",x"49",x"c7"),
   231 => (x"ff",x"b7",x"a9",x"06"),
   232 => (x"c3",x"d6",x"87",x"c8"),
   233 => (x"c0",x"1e",x"c8",x"66"),
   234 => (x"4a",x"75",x"82",x"72"),
   235 => (x"1e",x"27",x"15",x"15"),
   236 => (x"00",x"00",x"0f",x"c8"),
   237 => (x"86",x"70",x"4a",x"c8"),
   238 => (x"a6",x"49",x"72",x"79"),
   239 => (x"76",x"49",x"24",x"79"),
   240 => (x"c8",x"c0",x"85",x"c8"),
   241 => (x"c0",x"8b",x"c8",x"66"),
   242 => (x"49",x"6e",x"b7",x"a9"),
   243 => (x"02",x"c1",x"de",x"87"),
   244 => (x"27",x"60",x"18",x"00"),
   245 => (x"00",x"bf",x"1e",x"75"),
   246 => (x"1e",x"27",x"af",x"02"),
   247 => (x"00",x"00",x"0f",x"c8"),
   248 => (x"86",x"27",x"68",x"18"),
   249 => (x"00",x"00",x"49",x"c0"),
   250 => (x"e0",x"51",x"27",x"69"),
   251 => (x"18",x"00",x"00",x"bf"),
   252 => (x"1e",x"cc",x"66",x"1e"),
   253 => (x"27",x"af",x"02",x"00"),
   254 => (x"00",x"0f",x"c8",x"86"),
   255 => (x"27",x"71",x"18",x"00"),
   256 => (x"00",x"49",x"c0",x"e0"),
   257 => (x"51",x"27",x"72",x"18"),
   258 => (x"00",x"00",x"bf",x"1e"),
   259 => (x"c4",x"66",x"1e",x"27"),
   260 => (x"af",x"02",x"00",x"00"),
   261 => (x"0f",x"c8",x"86",x"27"),
   262 => (x"7a",x"18",x"00",x"00"),
   263 => (x"49",x"c0",x"51",x"27"),
   264 => (x"60",x"18",x"00",x"00"),
   265 => (x"bf",x"1e",x"27",x"9e"),
   266 => (x"0d",x"00",x"00",x"0f"),
   267 => (x"c4",x"86",x"73",x"49"),
   268 => (x"c7",x"ff",x"b7",x"a9"),
   269 => (x"01",x"fd",x"eb",x"87"),
   270 => (x"c0",x"fe",x"87",x"27"),
   271 => (x"c2",x"15",x"00",x"00"),
   272 => (x"1e",x"27",x"9e",x"0d"),
   273 => (x"00",x"00",x"0f",x"c4"),
   274 => (x"86",x"c0",x"ed",x"87"),
   275 => (x"27",x"d7",x"15",x"00"),
   276 => (x"00",x"1e",x"27",x"9e"),
   277 => (x"0d",x"00",x"00",x"0f"),
   278 => (x"c4",x"86",x"27",x"f3"),
   279 => (x"15",x"00",x"00",x"1e"),
   280 => (x"27",x"b5",x"14",x"00"),
   281 => (x"00",x"0f",x"c4",x"86"),
   282 => (x"c0",x"ce",x"87",x"27"),
   283 => (x"52",x"16",x"00",x"00"),
   284 => (x"1e",x"27",x"9e",x"0d"),
   285 => (x"00",x"00",x"0f",x"c4"),
   286 => (x"86",x"ff",x"fd",x"87"),
   287 => (x"cc",x"86",x"26",x"4d"),
   288 => (x"26",x"4c",x"26",x"4b"),
   289 => (x"26",x"4a",x"26",x"4f"),
   290 => (x"0e",x"5e",x"5a",x"5b"),
   291 => (x"5c",x"5d",x"0e",x"d4"),
   292 => (x"66",x"4d",x"c0",x"4c"),
   293 => (x"dc",x"66",x"49",x"c0"),
   294 => (x"b7",x"a9",x"06",x"c0"),
   295 => (x"f2",x"87",x"15",x"4b"),
   296 => (x"d8",x"33",x"b7",x"2b"),
   297 => (x"d8",x"a6",x"bf",x"97"),
   298 => (x"bf",x"4a",x"d8",x"32"),
   299 => (x"b7",x"2a",x"d8",x"66"),
   300 => (x"48",x"c1",x"80",x"dc"),
   301 => (x"a6",x"58",x"73",x"49"),
   302 => (x"72",x"b7",x"a9",x"02"),
   303 => (x"c0",x"c5",x"87",x"c1"),
   304 => (x"48",x"c0",x"ce",x"87"),
   305 => (x"c1",x"84",x"74",x"49"),
   306 => (x"dc",x"66",x"b7",x"a9"),
   307 => (x"04",x"ff",x"ce",x"87"),
   308 => (x"c0",x"48",x"26",x"4d"),
   309 => (x"26",x"4c",x"26",x"4b"),
   310 => (x"26",x"4a",x"26",x"4f"),
   311 => (x"0e",x"5e",x"5a",x"5b"),
   312 => (x"5c",x"5d",x"0e",x"27"),
   313 => (x"b4",x"1a",x"00",x"00"),
   314 => (x"49",x"ff",x"79",x"27"),
   315 => (x"c4",x"1a",x"00",x"00"),
   316 => (x"49",x"c0",x"79",x"27"),
   317 => (x"62",x"17",x"00",x"00"),
   318 => (x"1e",x"27",x"b5",x"14"),
   319 => (x"00",x"00",x"0f",x"c4"),
   320 => (x"86",x"27",x"b0",x"18"),
   321 => (x"00",x"00",x"bf",x"1e"),
   322 => (x"c0",x"1e",x"27",x"9f"),
   323 => (x"13",x"00",x"00",x"0f"),
   324 => (x"c8",x"86",x"70",x"4a"),
   325 => (x"72",x"9a",x"05",x"c0"),
   326 => (x"d3",x"87",x"27",x"70"),
   327 => (x"16",x"00",x"00",x"1e"),
   328 => (x"27",x"b5",x"14",x"00"),
   329 => (x"00",x"0f",x"c4",x"86"),
   330 => (x"c0",x"48",x"cf",x"ed"),
   331 => (x"87",x"27",x"6f",x"17"),
   332 => (x"00",x"00",x"1e",x"27"),
   333 => (x"b5",x"14",x"00",x"00"),
   334 => (x"0f",x"c4",x"86",x"c0"),
   335 => (x"4c",x"27",x"a0",x"18"),
   336 => (x"00",x"00",x"49",x"c1"),
   337 => (x"79",x"c8",x"1e",x"27"),
   338 => (x"86",x"17",x"00",x"00"),
   339 => (x"1e",x"27",x"e6",x"18"),
   340 => (x"00",x"00",x"bf",x"1e"),
   341 => (x"27",x"88",x"04",x"00"),
   342 => (x"00",x"0f",x"cc",x"86"),
   343 => (x"70",x"4a",x"72",x"9a"),
   344 => (x"05",x"c0",x"c8",x"87"),
   345 => (x"27",x"a0",x"18",x"00"),
   346 => (x"00",x"49",x"c0",x"79"),
   347 => (x"c8",x"1e",x"27",x"8f"),
   348 => (x"17",x"00",x"00",x"1e"),
   349 => (x"27",x"02",x"19",x"00"),
   350 => (x"00",x"bf",x"1e",x"27"),
   351 => (x"88",x"04",x"00",x"00"),
   352 => (x"0f",x"cc",x"86",x"70"),
   353 => (x"4a",x"72",x"9a",x"05"),
   354 => (x"c0",x"c8",x"87",x"27"),
   355 => (x"a0",x"18",x"00",x"00"),
   356 => (x"49",x"c0",x"79",x"c8"),
   357 => (x"1e",x"27",x"98",x"17"),
   358 => (x"00",x"00",x"1e",x"27"),
   359 => (x"02",x"19",x"00",x"00"),
   360 => (x"bf",x"1e",x"27",x"88"),
   361 => (x"04",x"00",x"00",x"0f"),
   362 => (x"cc",x"86",x"70",x"4a"),
   363 => (x"72",x"9a",x"05",x"c0"),
   364 => (x"d3",x"87",x"27",x"84"),
   365 => (x"16",x"00",x"00",x"1e"),
   366 => (x"27",x"b5",x"14",x"00"),
   367 => (x"00",x"0f",x"c4",x"86"),
   368 => (x"c0",x"48",x"cd",x"d5"),
   369 => (x"87",x"27",x"a0",x"18"),
   370 => (x"00",x"00",x"bf",x"1e"),
   371 => (x"27",x"a1",x"17",x"00"),
   372 => (x"00",x"1e",x"27",x"d9"),
   373 => (x"00",x"00",x"00",x"0f"),
   374 => (x"c8",x"86",x"27",x"a0"),
   375 => (x"18",x"00",x"00",x"bf"),
   376 => (x"02",x"c2",x"d6",x"87"),
   377 => (x"27",x"b0",x"18",x"00"),
   378 => (x"00",x"4b",x"27",x"78"),
   379 => (x"1a",x"00",x"00",x"bf"),
   380 => (x"4c",x"27",x"b0",x"1a"),
   381 => (x"00",x"00",x"9f",x"bf"),
   382 => (x"4a",x"72",x"49",x"c5"),
   383 => (x"d6",x"ea",x"b7",x"a9"),
   384 => (x"05",x"c0",x"d4",x"87"),
   385 => (x"73",x"4a",x"c7",x"c8"),
   386 => (x"82",x"6a",x"1e",x"27"),
   387 => (x"25",x"02",x"00",x"00"),
   388 => (x"0f",x"c4",x"86",x"70"),
   389 => (x"4c",x"c0",x"e6",x"87"),
   390 => (x"73",x"4a",x"c8",x"c0"),
   391 => (x"82",x"9f",x"6a",x"4a"),
   392 => (x"72",x"49",x"ca",x"e9"),
   393 => (x"d5",x"b7",x"a9",x"02"),
   394 => (x"c0",x"d3",x"87",x"27"),
   395 => (x"bb",x"16",x"00",x"00"),
   396 => (x"1e",x"27",x"b5",x"14"),
   397 => (x"00",x"00",x"0f",x"c4"),
   398 => (x"86",x"c0",x"48",x"cb"),
   399 => (x"dc",x"87",x"74",x"1e"),
   400 => (x"27",x"d9",x"16",x"00"),
   401 => (x"00",x"1e",x"27",x"d9"),
   402 => (x"00",x"00",x"00",x"0f"),
   403 => (x"c8",x"86",x"27",x"b0"),
   404 => (x"18",x"00",x"00",x"bf"),
   405 => (x"1e",x"74",x"1e",x"27"),
   406 => (x"9f",x"13",x"00",x"00"),
   407 => (x"0f",x"c8",x"86",x"70"),
   408 => (x"4a",x"72",x"9a",x"05"),
   409 => (x"c0",x"c5",x"87",x"c0"),
   410 => (x"48",x"ca",x"ee",x"87"),
   411 => (x"27",x"f1",x"16",x"00"),
   412 => (x"00",x"1e",x"27",x"b5"),
   413 => (x"14",x"00",x"00",x"0f"),
   414 => (x"c4",x"86",x"27",x"b4"),
   415 => (x"17",x"00",x"00",x"1e"),
   416 => (x"27",x"d9",x"00",x"00"),
   417 => (x"00",x"0f",x"c4",x"86"),
   418 => (x"c8",x"1e",x"27",x"cc"),
   419 => (x"17",x"00",x"00",x"1e"),
   420 => (x"27",x"02",x"19",x"00"),
   421 => (x"00",x"bf",x"1e",x"27"),
   422 => (x"88",x"04",x"00",x"00"),
   423 => (x"0f",x"cc",x"86",x"70"),
   424 => (x"4a",x"72",x"9a",x"05"),
   425 => (x"c0",x"cb",x"87",x"27"),
   426 => (x"c4",x"1a",x"00",x"00"),
   427 => (x"49",x"c1",x"79",x"c1"),
   428 => (x"c0",x"87",x"c8",x"1e"),
   429 => (x"27",x"d5",x"17",x"00"),
   430 => (x"00",x"1e",x"27",x"e6"),
   431 => (x"18",x"00",x"00",x"bf"),
   432 => (x"1e",x"27",x"88",x"04"),
   433 => (x"00",x"00",x"0f",x"cc"),
   434 => (x"86",x"70",x"4a",x"72"),
   435 => (x"9a",x"02",x"c0",x"e1"),
   436 => (x"87",x"27",x"18",x"17"),
   437 => (x"00",x"00",x"1e",x"27"),
   438 => (x"d9",x"00",x"00",x"00"),
   439 => (x"0f",x"c4",x"86",x"27"),
   440 => (x"35",x"17",x"00",x"00"),
   441 => (x"1e",x"27",x"b5",x"14"),
   442 => (x"00",x"00",x"0f",x"c4"),
   443 => (x"86",x"c0",x"48",x"c8"),
   444 => (x"e8",x"87",x"27",x"ae"),
   445 => (x"1a",x"00",x"00",x"97"),
   446 => (x"bf",x"4a",x"72",x"49"),
   447 => (x"c1",x"d5",x"b7",x"a9"),
   448 => (x"05",x"c0",x"d2",x"87"),
   449 => (x"27",x"af",x"1a",x"00"),
   450 => (x"00",x"97",x"bf",x"4a"),
   451 => (x"72",x"49",x"c2",x"ea"),
   452 => (x"b7",x"a9",x"02",x"c0"),
   453 => (x"c5",x"87",x"c0",x"48"),
   454 => (x"c7",x"ff",x"87",x"27"),
   455 => (x"b0",x"18",x"00",x"00"),
   456 => (x"97",x"bf",x"4a",x"72"),
   457 => (x"49",x"c3",x"e9",x"b7"),
   458 => (x"a9",x"02",x"c0",x"d7"),
   459 => (x"87",x"27",x"b0",x"18"),
   460 => (x"00",x"00",x"97",x"bf"),
   461 => (x"4a",x"72",x"49",x"c3"),
   462 => (x"eb",x"b7",x"a9",x"02"),
   463 => (x"c0",x"c5",x"87",x"c0"),
   464 => (x"48",x"c7",x"d6",x"87"),
   465 => (x"27",x"bb",x"18",x"00"),
   466 => (x"00",x"97",x"bf",x"4a"),
   467 => (x"72",x"9a",x"05",x"c0"),
   468 => (x"d1",x"87",x"27",x"bc"),
   469 => (x"18",x"00",x"00",x"97"),
   470 => (x"bf",x"4a",x"72",x"49"),
   471 => (x"c2",x"b7",x"a9",x"02"),
   472 => (x"c0",x"c5",x"87",x"c0"),
   473 => (x"48",x"c6",x"f2",x"87"),
   474 => (x"27",x"bd",x"18",x"00"),
   475 => (x"00",x"97",x"bf",x"48"),
   476 => (x"27",x"9c",x"18",x"00"),
   477 => (x"00",x"58",x"27",x"9c"),
   478 => (x"18",x"00",x"00",x"bf"),
   479 => (x"48",x"c1",x"88",x"27"),
   480 => (x"d8",x"1a",x"00",x"00"),
   481 => (x"58",x"27",x"be",x"18"),
   482 => (x"00",x"00",x"97",x"bf"),
   483 => (x"4a",x"74",x"82",x"27"),
   484 => (x"bf",x"18",x"00",x"00"),
   485 => (x"97",x"bf",x"4b",x"c8"),
   486 => (x"33",x"73",x"48",x"72"),
   487 => (x"80",x"27",x"a4",x"18"),
   488 => (x"00",x"00",x"58",x"27"),
   489 => (x"c0",x"18",x"00",x"00"),
   490 => (x"97",x"bf",x"48",x"27"),
   491 => (x"cc",x"1a",x"00",x"00"),
   492 => (x"58",x"27",x"c4",x"1a"),
   493 => (x"00",x"00",x"bf",x"02"),
   494 => (x"c3",x"e5",x"87",x"c8"),
   495 => (x"1e",x"27",x"59",x"17"),
   496 => (x"00",x"00",x"1e",x"27"),
   497 => (x"02",x"19",x"00",x"00"),
   498 => (x"bf",x"1e",x"27",x"88"),
   499 => (x"04",x"00",x"00",x"0f"),
   500 => (x"cc",x"86",x"70",x"4a"),
   501 => (x"72",x"9a",x"02",x"c0"),
   502 => (x"c5",x"87",x"c0",x"48"),
   503 => (x"c4",x"fb",x"87",x"27"),
   504 => (x"9c",x"18",x"00",x"00"),
   505 => (x"bf",x"48",x"c4",x"30"),
   506 => (x"27",x"d0",x"1a",x"00"),
   507 => (x"00",x"58",x"27",x"9c"),
   508 => (x"18",x"00",x"00",x"bf"),
   509 => (x"4b",x"27",x"d4",x"1a"),
   510 => (x"00",x"00",x"49",x"73"),
   511 => (x"79",x"27",x"d5",x"18"),
   512 => (x"00",x"00",x"97",x"bf"),
   513 => (x"4a",x"c8",x"32",x"27"),
   514 => (x"d4",x"18",x"00",x"00"),
   515 => (x"97",x"bf",x"4c",x"72"),
   516 => (x"4a",x"74",x"82",x"27"),
   517 => (x"d6",x"18",x"00",x"00"),
   518 => (x"97",x"bf",x"4c",x"d0"),
   519 => (x"34",x"72",x"4a",x"74"),
   520 => (x"82",x"27",x"d7",x"18"),
   521 => (x"00",x"00",x"97",x"bf"),
   522 => (x"4c",x"d8",x"34",x"72"),
   523 => (x"4a",x"74",x"82",x"27"),
   524 => (x"dc",x"1a",x"00",x"00"),
   525 => (x"49",x"72",x"79",x"72"),
   526 => (x"4a",x"27",x"cc",x"1a"),
   527 => (x"00",x"00",x"bf",x"92"),
   528 => (x"72",x"4a",x"27",x"a4"),
   529 => (x"18",x"00",x"00",x"bf"),
   530 => (x"82",x"27",x"c0",x"1a"),
   531 => (x"00",x"00",x"49",x"72"),
   532 => (x"79",x"27",x"dd",x"18"),
   533 => (x"00",x"00",x"97",x"bf"),
   534 => (x"4c",x"c8",x"34",x"27"),
   535 => (x"dc",x"18",x"00",x"00"),
   536 => (x"97",x"bf",x"4d",x"74"),
   537 => (x"4c",x"75",x"84",x"27"),
   538 => (x"de",x"18",x"00",x"00"),
   539 => (x"97",x"bf",x"4d",x"d0"),
   540 => (x"35",x"74",x"4c",x"75"),
   541 => (x"84",x"27",x"df",x"18"),
   542 => (x"00",x"00",x"97",x"bf"),
   543 => (x"4d",x"cf",x"9d",x"d8"),
   544 => (x"35",x"74",x"4c",x"75"),
   545 => (x"84",x"27",x"b0",x"1a"),
   546 => (x"00",x"00",x"49",x"74"),
   547 => (x"79",x"c2",x"8c",x"73"),
   548 => (x"4b",x"74",x"93",x"73"),
   549 => (x"48",x"72",x"80",x"27"),
   550 => (x"bc",x"1a",x"00",x"00"),
   551 => (x"58",x"c1",x"f8",x"87"),
   552 => (x"27",x"c2",x"18",x"00"),
   553 => (x"00",x"97",x"bf",x"4a"),
   554 => (x"c8",x"32",x"27",x"c1"),
   555 => (x"18",x"00",x"00",x"97"),
   556 => (x"bf",x"4b",x"72",x"4a"),
   557 => (x"73",x"82",x"27",x"d0"),
   558 => (x"1a",x"00",x"00",x"49"),
   559 => (x"72",x"79",x"c5",x"32"),
   560 => (x"c7",x"ff",x"82",x"c9"),
   561 => (x"b7",x"2a",x"27",x"d4"),
   562 => (x"1a",x"00",x"00",x"49"),
   563 => (x"72",x"79",x"27",x"c7"),
   564 => (x"18",x"00",x"00",x"97"),
   565 => (x"bf",x"4b",x"c8",x"33"),
   566 => (x"27",x"c6",x"18",x"00"),
   567 => (x"00",x"97",x"bf",x"4c"),
   568 => (x"73",x"4b",x"74",x"83"),
   569 => (x"27",x"dc",x"1a",x"00"),
   570 => (x"00",x"49",x"73",x"79"),
   571 => (x"73",x"4b",x"27",x"cc"),
   572 => (x"1a",x"00",x"00",x"bf"),
   573 => (x"93",x"73",x"4b",x"27"),
   574 => (x"a4",x"18",x"00",x"00"),
   575 => (x"bf",x"83",x"27",x"bc"),
   576 => (x"1a",x"00",x"00",x"49"),
   577 => (x"73",x"79",x"27",x"b0"),
   578 => (x"1a",x"00",x"00",x"49"),
   579 => (x"c0",x"79",x"73",x"48"),
   580 => (x"72",x"80",x"27",x"c0"),
   581 => (x"1a",x"00",x"00",x"58"),
   582 => (x"c1",x"48",x"26",x"4d"),
   583 => (x"26",x"4c",x"26",x"4b"),
   584 => (x"26",x"4a",x"26",x"4f"),
   585 => (x"0e",x"5e",x"5a",x"5b"),
   586 => (x"5c",x"5d",x"0e",x"27"),
   587 => (x"c4",x"1a",x"00",x"00"),
   588 => (x"bf",x"02",x"c0",x"cf"),
   589 => (x"87",x"d4",x"66",x"4b"),
   590 => (x"c7",x"b7",x"2b",x"d4"),
   591 => (x"66",x"4c",x"c1",x"ff"),
   592 => (x"9c",x"c0",x"cc",x"87"),
   593 => (x"d4",x"66",x"4b",x"c8"),
   594 => (x"b7",x"2b",x"d4",x"66"),
   595 => (x"4c",x"c3",x"ff",x"9c"),
   596 => (x"73",x"49",x"27",x"b4"),
   597 => (x"1a",x"00",x"00",x"bf"),
   598 => (x"a9",x"02",x"c0",x"ef"),
   599 => (x"87",x"27",x"b0",x"18"),
   600 => (x"00",x"00",x"bf",x"1e"),
   601 => (x"27",x"a4",x"18",x"00"),
   602 => (x"00",x"bf",x"4a",x"73"),
   603 => (x"82",x"72",x"1e",x"27"),
   604 => (x"9f",x"13",x"00",x"00"),
   605 => (x"0f",x"c8",x"86",x"70"),
   606 => (x"4a",x"72",x"9a",x"05"),
   607 => (x"c0",x"c5",x"87",x"c0"),
   608 => (x"48",x"c1",x"d4",x"87"),
   609 => (x"27",x"b4",x"1a",x"00"),
   610 => (x"00",x"49",x"73",x"79"),
   611 => (x"27",x"c4",x"1a",x"00"),
   612 => (x"00",x"bf",x"02",x"c0"),
   613 => (x"e4",x"87",x"74",x"4a"),
   614 => (x"c4",x"92",x"72",x"4a"),
   615 => (x"27",x"b0",x"18",x"00"),
   616 => (x"00",x"bf",x"82",x"6a"),
   617 => (x"1e",x"27",x"25",x"02"),
   618 => (x"00",x"00",x"0f",x"c4"),
   619 => (x"86",x"70",x"4a",x"72"),
   620 => (x"4d",x"cf",x"ff",x"ff"),
   621 => (x"ff",x"ff",x"9d",x"c0"),
   622 => (x"dc",x"87",x"74",x"4a"),
   623 => (x"c2",x"92",x"72",x"4a"),
   624 => (x"27",x"b0",x"18",x"00"),
   625 => (x"00",x"bf",x"82",x"9f"),
   626 => (x"6a",x"4a",x"72",x"1e"),
   627 => (x"27",x"67",x"02",x"00"),
   628 => (x"00",x"0f",x"c4",x"86"),
   629 => (x"70",x"4d",x"75",x"48"),
   630 => (x"26",x"4d",x"26",x"4c"),
   631 => (x"26",x"4b",x"26",x"4a"),
   632 => (x"26",x"4f",x"0e",x"5e"),
   633 => (x"5a",x"5b",x"5c",x"5d"),
   634 => (x"0e",x"d0",x"8e",x"cf"),
   635 => (x"ff",x"ff",x"ff",x"f8"),
   636 => (x"4d",x"c0",x"4c",x"27"),
   637 => (x"b4",x"1a",x"00",x"00"),
   638 => (x"49",x"ff",x"79",x"76"),
   639 => (x"49",x"27",x"b0",x"1a"),
   640 => (x"00",x"00",x"bf",x"79"),
   641 => (x"27",x"bc",x"1a",x"00"),
   642 => (x"00",x"bf",x"4b",x"27"),
   643 => (x"c4",x"1a",x"00",x"00"),
   644 => (x"bf",x"02",x"c0",x"cc"),
   645 => (x"87",x"27",x"9c",x"18"),
   646 => (x"00",x"00",x"bf",x"4a"),
   647 => (x"c4",x"32",x"c0",x"c9"),
   648 => (x"87",x"27",x"d4",x"1a"),
   649 => (x"00",x"00",x"bf",x"4a"),
   650 => (x"c4",x"32",x"c8",x"a6"),
   651 => (x"49",x"72",x"79",x"c4"),
   652 => (x"a6",x"49",x"73",x"79"),
   653 => (x"c0",x"4b",x"c8",x"66"),
   654 => (x"49",x"c0",x"a9",x"06"),
   655 => (x"c4",x"dd",x"87",x"73"),
   656 => (x"4a",x"cf",x"9a",x"72"),
   657 => (x"9a",x"05",x"c0",x"f4"),
   658 => (x"87",x"c4",x"66",x"1e"),
   659 => (x"27",x"c5",x"0b",x"00"),
   660 => (x"00",x"1e",x"27",x"d9"),
   661 => (x"00",x"00",x"00",x"0f"),
   662 => (x"c8",x"86",x"27",x"b0"),
   663 => (x"18",x"00",x"00",x"bf"),
   664 => (x"1e",x"c8",x"66",x"1e"),
   665 => (x"cc",x"66",x"48",x"c1"),
   666 => (x"80",x"d0",x"a6",x"58"),
   667 => (x"27",x"9f",x"13",x"00"),
   668 => (x"00",x"0f",x"c8",x"86"),
   669 => (x"27",x"b0",x"18",x"00"),
   670 => (x"00",x"4c",x"c0",x"c3"),
   671 => (x"87",x"c0",x"e0",x"84"),
   672 => (x"97",x"6c",x"4a",x"cc"),
   673 => (x"a6",x"49",x"73",x"79"),
   674 => (x"72",x"9a",x"02",x"c3"),
   675 => (x"c3",x"87",x"97",x"6c"),
   676 => (x"4a",x"cc",x"a6",x"49"),
   677 => (x"73",x"79",x"72",x"49"),
   678 => (x"c3",x"e5",x"b7",x"a9"),
   679 => (x"02",x"c2",x"f1",x"87"),
   680 => (x"74",x"4a",x"cb",x"82"),
   681 => (x"97",x"6a",x"4a",x"d8"),
   682 => (x"9a",x"cc",x"a6",x"49"),
   683 => (x"73",x"79",x"72",x"9a"),
   684 => (x"05",x"c2",x"dd",x"87"),
   685 => (x"cb",x"1e",x"c0",x"ec"),
   686 => (x"66",x"1e",x"74",x"1e"),
   687 => (x"27",x"88",x"04",x"00"),
   688 => (x"00",x"0f",x"cc",x"86"),
   689 => (x"70",x"4a",x"cc",x"a6"),
   690 => (x"49",x"73",x"79",x"72"),
   691 => (x"9a",x"05",x"c2",x"c0"),
   692 => (x"87",x"74",x"4a",x"dc"),
   693 => (x"82",x"6a",x"1e",x"27"),
   694 => (x"25",x"02",x"00",x"00"),
   695 => (x"0f",x"c4",x"86",x"70"),
   696 => (x"4b",x"c0",x"e4",x"66"),
   697 => (x"4a",x"c4",x"82",x"73"),
   698 => (x"7a",x"74",x"4a",x"da"),
   699 => (x"82",x"9f",x"6a",x"4a"),
   700 => (x"72",x"1e",x"27",x"67"),
   701 => (x"02",x"00",x"00",x"0f"),
   702 => (x"c4",x"86",x"c4",x"a6"),
   703 => (x"58",x"27",x"c4",x"1a"),
   704 => (x"00",x"00",x"bf",x"02"),
   705 => (x"c0",x"de",x"87",x"74"),
   706 => (x"4a",x"d4",x"82",x"9f"),
   707 => (x"6a",x"4a",x"72",x"1e"),
   708 => (x"27",x"67",x"02",x"00"),
   709 => (x"00",x"0f",x"c4",x"86"),
   710 => (x"70",x"4a",x"c0",x"ff"),
   711 => (x"ff",x"9a",x"72",x"4d"),
   712 => (x"d0",x"35",x"c0",x"c2"),
   713 => (x"87",x"c0",x"4d",x"75"),
   714 => (x"4b",x"6e",x"83",x"c0"),
   715 => (x"e4",x"66",x"4a",x"c8"),
   716 => (x"82",x"73",x"7a",x"c0"),
   717 => (x"e4",x"a6",x"bf",x"49"),
   718 => (x"c0",x"79",x"c0",x"e8"),
   719 => (x"66",x"1e",x"27",x"e2"),
   720 => (x"0b",x"00",x"00",x"1e"),
   721 => (x"27",x"d9",x"00",x"00"),
   722 => (x"00",x"0f",x"c8",x"86"),
   723 => (x"c1",x"48",x"c1",x"e2"),
   724 => (x"87",x"c1",x"83",x"73"),
   725 => (x"49",x"c8",x"66",x"a9"),
   726 => (x"04",x"fb",x"e3",x"87"),
   727 => (x"cf",x"ff",x"ff",x"ff"),
   728 => (x"f8",x"4d",x"27",x"c4"),
   729 => (x"1a",x"00",x"00",x"bf"),
   730 => (x"02",x"c1",x"c5",x"87"),
   731 => (x"6e",x"1e",x"27",x"24"),
   732 => (x"09",x"00",x"00",x"0f"),
   733 => (x"c4",x"86",x"c4",x"a6"),
   734 => (x"58",x"6e",x"1e",x"27"),
   735 => (x"f3",x"0b",x"00",x"00"),
   736 => (x"1e",x"27",x"d9",x"00"),
   737 => (x"00",x"00",x"0f",x"c8"),
   738 => (x"86",x"6e",x"4a",x"75"),
   739 => (x"9a",x"72",x"49",x"75"),
   740 => (x"a9",x"02",x"c0",x"dc"),
   741 => (x"87",x"6e",x"4a",x"c2"),
   742 => (x"8a",x"72",x"4a",x"27"),
   743 => (x"9c",x"18",x"00",x"00"),
   744 => (x"bf",x"92",x"27",x"c0"),
   745 => (x"1a",x"00",x"00",x"bf"),
   746 => (x"48",x"72",x"80",x"c8"),
   747 => (x"a6",x"58",x"fa",x"c3"),
   748 => (x"87",x"c0",x"48",x"cf"),
   749 => (x"ff",x"ff",x"ff",x"f8"),
   750 => (x"4d",x"d0",x"86",x"26"),
   751 => (x"4d",x"26",x"4c",x"26"),
   752 => (x"4b",x"26",x"4a",x"26"),
   753 => (x"4f",x"52",x"65",x"61"),
   754 => (x"64",x"69",x"6e",x"67"),
   755 => (x"20",x"64",x"69",x"72"),
   756 => (x"65",x"63",x"74",x"6f"),
   757 => (x"72",x"79",x"20",x"73"),
   758 => (x"65",x"63",x"74",x"6f"),
   759 => (x"72",x"20",x"25",x"64"),
   760 => (x"0a",x"00",x"66",x"69"),
   761 => (x"6c",x"65",x"20",x"22"),
   762 => (x"25",x"73",x"22",x"20"),
   763 => (x"66",x"6f",x"75",x"6e"),
   764 => (x"64",x"0d",x"00",x"47"),
   765 => (x"65",x"74",x"46",x"41"),
   766 => (x"54",x"4c",x"69",x"6e"),
   767 => (x"6b",x"20",x"72",x"65"),
   768 => (x"74",x"75",x"72",x"6e"),
   769 => (x"65",x"64",x"20",x"25"),
   770 => (x"64",x"0a",x"00",x"0e"),
   771 => (x"5e",x"5a",x"5b",x"5c"),
   772 => (x"5d",x"0e",x"1e",x"d8"),
   773 => (x"66",x"1e",x"27",x"90"),
   774 => (x"18",x"00",x"00",x"bf"),
   775 => (x"1e",x"27",x"e2",x"09"),
   776 => (x"00",x"00",x"0f",x"c8"),
   777 => (x"86",x"70",x"4a",x"72"),
   778 => (x"9a",x"02",x"c2",x"e0"),
   779 => (x"87",x"27",x"94",x"18"),
   780 => (x"00",x"00",x"bf",x"4a"),
   781 => (x"c7",x"ff",x"82",x"c9"),
   782 => (x"b7",x"2a",x"76",x"49"),
   783 => (x"72",x"79",x"c0",x"4d"),
   784 => (x"c0",x"4c",x"6e",x"49"),
   785 => (x"c0",x"b7",x"a9",x"06"),
   786 => (x"c2",x"d8",x"87",x"27"),
   787 => (x"c0",x"1a",x"00",x"00"),
   788 => (x"bf",x"4a",x"27",x"98"),
   789 => (x"18",x"00",x"00",x"bf"),
   790 => (x"4b",x"c2",x"8b",x"73"),
   791 => (x"4b",x"27",x"9c",x"18"),
   792 => (x"00",x"00",x"bf",x"93"),
   793 => (x"72",x"4a",x"73",x"82"),
   794 => (x"27",x"d8",x"1a",x"00"),
   795 => (x"00",x"bf",x"4b",x"74"),
   796 => (x"9b",x"72",x"4a",x"73"),
   797 => (x"82",x"dc",x"66",x"1e"),
   798 => (x"72",x"1e",x"27",x"9f"),
   799 => (x"13",x"00",x"00",x"0f"),
   800 => (x"c8",x"86",x"70",x"4a"),
   801 => (x"72",x"9a",x"05",x"c0"),
   802 => (x"c5",x"87",x"c0",x"48"),
   803 => (x"c1",x"db",x"87",x"c1"),
   804 => (x"84",x"27",x"d8",x"1a"),
   805 => (x"00",x"00",x"bf",x"4a"),
   806 => (x"74",x"9a",x"72",x"9a"),
   807 => (x"05",x"c0",x"d5",x"87"),
   808 => (x"27",x"98",x"18",x"00"),
   809 => (x"00",x"bf",x"1e",x"27"),
   810 => (x"24",x"09",x"00",x"00"),
   811 => (x"0f",x"c4",x"86",x"27"),
   812 => (x"98",x"18",x"00",x"00"),
   813 => (x"58",x"dc",x"66",x"48"),
   814 => (x"c8",x"c0",x"80",x"c0"),
   815 => (x"e0",x"a6",x"58",x"c1"),
   816 => (x"85",x"75",x"49",x"6e"),
   817 => (x"b7",x"a9",x"04",x"fe"),
   818 => (x"c1",x"87",x"c0",x"d6"),
   819 => (x"87",x"d8",x"66",x"1e"),
   820 => (x"27",x"f5",x"0c",x"00"),
   821 => (x"00",x"1e",x"27",x"d9"),
   822 => (x"00",x"00",x"00",x"0f"),
   823 => (x"c8",x"86",x"c0",x"48"),
   824 => (x"c0",x"c7",x"87",x"27"),
   825 => (x"94",x"18",x"00",x"00"),
   826 => (x"bf",x"48",x"26",x"26"),
   827 => (x"4d",x"26",x"4c",x"26"),
   828 => (x"4b",x"26",x"4a",x"26"),
   829 => (x"4f",x"43",x"61",x"6e"),
   830 => (x"27",x"74",x"20",x"6f"),
   831 => (x"70",x"65",x"6e",x"20"),
   832 => (x"25",x"73",x"0a",x"00"),
   833 => (x"1e",x"72",x"1e",x"c8"),
   834 => (x"66",x"02",x"c0",x"d1"),
   835 => (x"87",x"27",x"80",x"18"),
   836 => (x"00",x"00",x"49",x"c8"),
   837 => (x"66",x"79",x"27",x"88"),
   838 => (x"18",x"00",x"00",x"49"),
   839 => (x"c0",x"79",x"27",x"88"),
   840 => (x"18",x"00",x"00",x"05"),
   841 => (x"c0",x"db",x"87",x"27"),
   842 => (x"80",x"18",x"00",x"00"),
   843 => (x"4a",x"72",x"48",x"c4"),
   844 => (x"80",x"27",x"80",x"18"),
   845 => (x"00",x"00",x"58",x"27"),
   846 => (x"84",x"18",x"00",x"00"),
   847 => (x"49",x"6a",x"79",x"c0"),
   848 => (x"ce",x"87",x"27",x"84"),
   849 => (x"18",x"00",x"00",x"48"),
   850 => (x"c8",x"30",x"27",x"84"),
   851 => (x"18",x"00",x"00",x"58"),
   852 => (x"27",x"88",x"18",x"00"),
   853 => (x"00",x"4a",x"c1",x"82"),
   854 => (x"72",x"48",x"c3",x"98"),
   855 => (x"27",x"88",x"18",x"00"),
   856 => (x"00",x"58",x"27",x"84"),
   857 => (x"18",x"00",x"00",x"4a"),
   858 => (x"d8",x"b7",x"2a",x"72"),
   859 => (x"48",x"26",x"4a",x"26"),
   860 => (x"4f",x"0e",x"5e",x"5a"),
   861 => (x"5b",x"0e",x"cc",x"66"),
   862 => (x"1e",x"fe",x"c8",x"87"),
   863 => (x"c4",x"86",x"70",x"4b"),
   864 => (x"c0",x"4a",x"73",x"9b"),
   865 => (x"02",x"c0",x"ce",x"87"),
   866 => (x"c1",x"82",x"c0",x"1e"),
   867 => (x"fd",x"f5",x"87",x"c4"),
   868 => (x"86",x"70",x"4b",x"ff"),
   869 => (x"ec",x"87",x"72",x"48"),
   870 => (x"26",x"4b",x"26",x"4a"),
   871 => (x"26",x"4f",x"0e",x"5e"),
   872 => (x"5a",x"5b",x"5c",x"5d"),
   873 => (x"0e",x"c8",x"8e",x"c0"),
   874 => (x"f6",x"e4",x"c0",x"c4"),
   875 => (x"4c",x"c0",x"f6",x"e4"),
   876 => (x"c0",x"c0",x"4b",x"dc"),
   877 => (x"66",x"1e",x"fe",x"f8"),
   878 => (x"87",x"c4",x"86",x"70"),
   879 => (x"4a",x"72",x"4d",x"c2"),
   880 => (x"85",x"76",x"49",x"c1"),
   881 => (x"79",x"d0",x"9f",x"7c"),
   882 => (x"c1",x"c0",x"c1",x"9f"),
   883 => (x"7b",x"9f",x"6b",x"4a"),
   884 => (x"c0",x"9f",x"7b",x"c0"),
   885 => (x"9f",x"7b",x"9f",x"6b"),
   886 => (x"48",x"c8",x"a6",x"58"),
   887 => (x"c4",x"c0",x"9a",x"72"),
   888 => (x"9a",x"02",x"c1",x"fe"),
   889 => (x"87",x"6e",x"02",x"c0"),
   890 => (x"e6",x"87",x"c4",x"66"),
   891 => (x"49",x"c8",x"c0",x"c6"),
   892 => (x"a9",x"05",x"c1",x"ee"),
   893 => (x"87",x"76",x"49",x"c0"),
   894 => (x"79",x"fa",x"eb",x"ca"),
   895 => (x"9f",x"7b",x"c1",x"9f"),
   896 => (x"7b",x"c0",x"9f",x"7b"),
   897 => (x"75",x"9f",x"7b",x"c0"),
   898 => (x"9f",x"7b",x"c0",x"9f"),
   899 => (x"7b",x"c1",x"d3",x"87"),
   900 => (x"75",x"4a",x"c1",x"b7"),
   901 => (x"2a",x"c8",x"c0",x"c0"),
   902 => (x"b2",x"c4",x"66",x"49"),
   903 => (x"72",x"a9",x"05",x"c1"),
   904 => (x"c1",x"87",x"dc",x"66"),
   905 => (x"1e",x"fb",x"dc",x"87"),
   906 => (x"c4",x"86",x"c4",x"a6"),
   907 => (x"58",x"75",x"4a",x"c1"),
   908 => (x"8d",x"72",x"9a",x"02"),
   909 => (x"c0",x"de",x"87",x"6e"),
   910 => (x"4c",x"74",x"97",x"7b"),
   911 => (x"74",x"9c",x"02",x"c0"),
   912 => (x"c9",x"87",x"c0",x"1e"),
   913 => (x"fa",x"fd",x"87",x"c4"),
   914 => (x"86",x"70",x"4c",x"75"),
   915 => (x"4a",x"c1",x"8d",x"72"),
   916 => (x"9a",x"05",x"ff",x"e4"),
   917 => (x"87",x"c0",x"f6",x"e4"),
   918 => (x"c0",x"c4",x"4c",x"d1"),
   919 => (x"9f",x"7c",x"c1",x"48"),
   920 => (x"c0",x"c6",x"87",x"d1"),
   921 => (x"9f",x"7c",x"fd",x"dc"),
   922 => (x"87",x"c8",x"86",x"26"),
   923 => (x"4d",x"26",x"4c",x"26"),
   924 => (x"4b",x"26",x"4a",x"26"),
   925 => (x"4f",x"0e",x"5e",x"5a"),
   926 => (x"5b",x"0e",x"dc",x"8e"),
   927 => (x"c0",x"f6",x"e4",x"c0"),
   928 => (x"c0",x"4b",x"ff",x"97"),
   929 => (x"7b",x"97",x"6b",x"48"),
   930 => (x"c4",x"a6",x"58",x"6e"),
   931 => (x"4a",x"c3",x"ff",x"9a"),
   932 => (x"ff",x"97",x"7b",x"c8"),
   933 => (x"32",x"97",x"6b",x"48"),
   934 => (x"c8",x"a6",x"58",x"c4"),
   935 => (x"66",x"48",x"c3",x"ff"),
   936 => (x"98",x"cc",x"a6",x"58"),
   937 => (x"72",x"4a",x"c8",x"66"),
   938 => (x"b2",x"ff",x"97",x"7b"),
   939 => (x"c8",x"32",x"97",x"6b"),
   940 => (x"48",x"d0",x"a6",x"58"),
   941 => (x"cc",x"66",x"48",x"c3"),
   942 => (x"ff",x"98",x"d4",x"a6"),
   943 => (x"58",x"72",x"4a",x"d0"),
   944 => (x"66",x"b2",x"ff",x"97"),
   945 => (x"7b",x"c8",x"32",x"13"),
   946 => (x"48",x"d8",x"a6",x"58"),
   947 => (x"d4",x"66",x"48",x"c3"),
   948 => (x"ff",x"98",x"dc",x"a6"),
   949 => (x"58",x"72",x"4a",x"d8"),
   950 => (x"66",x"b2",x"72",x"48"),
   951 => (x"dc",x"86",x"26",x"4b"),
   952 => (x"26",x"4a",x"26",x"4f"),
   953 => (x"0e",x"5e",x"5a",x"5b"),
   954 => (x"5c",x"5d",x"0e",x"1e"),
   955 => (x"c0",x"f6",x"e4",x"c0"),
   956 => (x"c0",x"4b",x"d8",x"66"),
   957 => (x"4a",x"c3",x"ff",x"9a"),
   958 => (x"72",x"97",x"7b",x"27"),
   959 => (x"e0",x"1a",x"00",x"00"),
   960 => (x"bf",x"05",x"c0",x"c9"),
   961 => (x"87",x"dc",x"66",x"48"),
   962 => (x"c9",x"30",x"c0",x"e0"),
   963 => (x"a6",x"58",x"dc",x"66"),
   964 => (x"4a",x"d8",x"b7",x"2a"),
   965 => (x"c3",x"ff",x"9a",x"72"),
   966 => (x"97",x"7b",x"dc",x"66"),
   967 => (x"4a",x"d0",x"b7",x"2a"),
   968 => (x"c3",x"ff",x"9a",x"72"),
   969 => (x"97",x"7b",x"dc",x"66"),
   970 => (x"4a",x"c8",x"b7",x"2a"),
   971 => (x"c3",x"ff",x"9a",x"72"),
   972 => (x"97",x"7b",x"dc",x"66"),
   973 => (x"4a",x"c3",x"ff",x"9a"),
   974 => (x"72",x"97",x"7b",x"d8"),
   975 => (x"66",x"4a",x"d0",x"b7"),
   976 => (x"2a",x"c3",x"ff",x"9a"),
   977 => (x"72",x"97",x"7b",x"97"),
   978 => (x"6b",x"48",x"c4",x"a6"),
   979 => (x"58",x"6e",x"4d",x"c3"),
   980 => (x"ff",x"9d",x"c9",x"f0"),
   981 => (x"ff",x"4c",x"75",x"49"),
   982 => (x"c3",x"ff",x"b7",x"a9"),
   983 => (x"05",x"c0",x"e1",x"87"),
   984 => (x"c3",x"ff",x"4a",x"ff"),
   985 => (x"97",x"7b",x"97",x"6b"),
   986 => (x"48",x"c4",x"a6",x"58"),
   987 => (x"6e",x"4d",x"72",x"9d"),
   988 => (x"c1",x"8c",x"74",x"9c"),
   989 => (x"02",x"c0",x"c9",x"87"),
   990 => (x"75",x"49",x"72",x"b7"),
   991 => (x"a9",x"02",x"ff",x"e2"),
   992 => (x"87",x"75",x"1e",x"27"),
   993 => (x"de",x"17",x"00",x"00"),
   994 => (x"1e",x"27",x"d9",x"00"),
   995 => (x"00",x"00",x"0f",x"c8"),
   996 => (x"86",x"75",x"48",x"26"),
   997 => (x"26",x"4d",x"26",x"4c"),
   998 => (x"26",x"4b",x"26",x"4a"),
   999 => (x"26",x"4f",x"0e",x"5e"),
  1000 => (x"5a",x"5b",x"0e",x"c0"),
  1001 => (x"f6",x"e4",x"c0",x"c0"),
  1002 => (x"4b",x"c0",x"4a",x"ff"),
  1003 => (x"97",x"7b",x"c1",x"82"),
  1004 => (x"72",x"49",x"c3",x"c8"),
  1005 => (x"b7",x"a9",x"04",x"ff"),
  1006 => (x"f1",x"87",x"26",x"4b"),
  1007 => (x"26",x"4a",x"26",x"4f"),
  1008 => (x"0e",x"5e",x"5a",x"5b"),
  1009 => (x"5c",x"5d",x"0e",x"c1"),
  1010 => (x"c0",x"c0",x"c0",x"c0"),
  1011 => (x"c0",x"4c",x"c0",x"f6"),
  1012 => (x"e4",x"c0",x"c0",x"4b"),
  1013 => (x"27",x"9e",x"0f",x"00"),
  1014 => (x"00",x"0f",x"c0",x"86"),
  1015 => (x"c4",x"f8",x"df",x"4d"),
  1016 => (x"c0",x"1e",x"c0",x"ff"),
  1017 => (x"f0",x"c1",x"f7",x"1e"),
  1018 => (x"27",x"e4",x"0e",x"00"),
  1019 => (x"00",x"0f",x"c8",x"86"),
  1020 => (x"70",x"4a",x"72",x"49"),
  1021 => (x"c1",x"b7",x"a9",x"05"),
  1022 => (x"c1",x"de",x"87",x"72"),
  1023 => (x"1e",x"27",x"87",x"10"),
  1024 => (x"00",x"00",x"1e",x"27"),
  1025 => (x"d9",x"00",x"00",x"00"),
  1026 => (x"0f",x"c8",x"86",x"ff"),
  1027 => (x"97",x"7b",x"74",x"1e"),
  1028 => (x"c0",x"e1",x"f0",x"c1"),
  1029 => (x"e9",x"1e",x"27",x"e4"),
  1030 => (x"0e",x"00",x"00",x"0f"),
  1031 => (x"c8",x"86",x"70",x"4a"),
  1032 => (x"72",x"9a",x"05",x"c0"),
  1033 => (x"d8",x"87",x"72",x"1e"),
  1034 => (x"27",x"7d",x"10",x"00"),
  1035 => (x"00",x"1e",x"27",x"d9"),
  1036 => (x"00",x"00",x"00",x"0f"),
  1037 => (x"c8",x"86",x"ff",x"97"),
  1038 => (x"7b",x"c1",x"48",x"c0"),
  1039 => (x"f5",x"87",x"72",x"1e"),
  1040 => (x"27",x"91",x"10",x"00"),
  1041 => (x"00",x"1e",x"27",x"d9"),
  1042 => (x"00",x"00",x"00",x"0f"),
  1043 => (x"c8",x"86",x"27",x"9e"),
  1044 => (x"0f",x"00",x"00",x"0f"),
  1045 => (x"c0",x"86",x"c0",x"d0"),
  1046 => (x"87",x"72",x"1e",x"27"),
  1047 => (x"9b",x"10",x"00",x"00"),
  1048 => (x"1e",x"27",x"d9",x"00"),
  1049 => (x"00",x"00",x"0f",x"c8"),
  1050 => (x"86",x"c1",x"8d",x"75"),
  1051 => (x"9d",x"05",x"fd",x"ef"),
  1052 => (x"87",x"c0",x"48",x"26"),
  1053 => (x"4d",x"26",x"4c",x"26"),
  1054 => (x"4b",x"26",x"4a",x"26"),
  1055 => (x"4f",x"43",x"4d",x"44"),
  1056 => (x"34",x"31",x"20",x"25"),
  1057 => (x"64",x"0a",x"00",x"43"),
  1058 => (x"4d",x"44",x"35",x"35"),
  1059 => (x"20",x"25",x"64",x"0a"),
  1060 => (x"00",x"43",x"4d",x"44"),
  1061 => (x"34",x"31",x"20",x"25"),
  1062 => (x"64",x"0a",x"00",x"43"),
  1063 => (x"4d",x"44",x"35",x"35"),
  1064 => (x"20",x"25",x"64",x"0a"),
  1065 => (x"00",x"0e",x"5e",x"5a"),
  1066 => (x"5b",x"5c",x"5d",x"0e"),
  1067 => (x"c0",x"ff",x"f0",x"c1"),
  1068 => (x"c1",x"4d",x"c0",x"f6"),
  1069 => (x"e4",x"c0",x"c0",x"4b"),
  1070 => (x"ff",x"97",x"7b",x"27"),
  1071 => (x"39",x"11",x"00",x"00"),
  1072 => (x"1e",x"27",x"b5",x"14"),
  1073 => (x"00",x"00",x"0f",x"c4"),
  1074 => (x"86",x"d3",x"4c",x"c0"),
  1075 => (x"1e",x"75",x"1e",x"27"),
  1076 => (x"e4",x"0e",x"00",x"00"),
  1077 => (x"0f",x"c8",x"86",x"70"),
  1078 => (x"4a",x"72",x"9a",x"05"),
  1079 => (x"c0",x"d8",x"87",x"72"),
  1080 => (x"1e",x"27",x"23",x"11"),
  1081 => (x"00",x"00",x"1e",x"27"),
  1082 => (x"d9",x"00",x"00",x"00"),
  1083 => (x"0f",x"c8",x"86",x"ff"),
  1084 => (x"97",x"7b",x"c1",x"48"),
  1085 => (x"c0",x"e2",x"87",x"72"),
  1086 => (x"1e",x"27",x"2e",x"11"),
  1087 => (x"00",x"00",x"1e",x"27"),
  1088 => (x"d9",x"00",x"00",x"00"),
  1089 => (x"0f",x"c8",x"86",x"27"),
  1090 => (x"9e",x"0f",x"00",x"00"),
  1091 => (x"0f",x"c0",x"86",x"c1"),
  1092 => (x"8c",x"74",x"9c",x"05"),
  1093 => (x"fe",x"f4",x"87",x"c0"),
  1094 => (x"48",x"26",x"4d",x"26"),
  1095 => (x"4c",x"26",x"4b",x"26"),
  1096 => (x"4a",x"26",x"4f",x"69"),
  1097 => (x"6e",x"69",x"74",x"20"),
  1098 => (x"25",x"64",x"0a",x"20"),
  1099 => (x"20",x"00",x"69",x"6e"),
  1100 => (x"69",x"74",x"20",x"25"),
  1101 => (x"64",x"0a",x"20",x"20"),
  1102 => (x"00",x"43",x"6d",x"64"),
  1103 => (x"5f",x"69",x"6e",x"69"),
  1104 => (x"74",x"0a",x"00",x"0e"),
  1105 => (x"5e",x"5a",x"5b",x"5c"),
  1106 => (x"5d",x"0e",x"1e",x"c0"),
  1107 => (x"f6",x"e4",x"c0",x"c0"),
  1108 => (x"4b",x"27",x"9e",x"0f"),
  1109 => (x"00",x"00",x"0f",x"c0"),
  1110 => (x"86",x"c6",x"ea",x"1e"),
  1111 => (x"c0",x"e1",x"f0",x"c1"),
  1112 => (x"c8",x"1e",x"27",x"e4"),
  1113 => (x"0e",x"00",x"00",x"0f"),
  1114 => (x"c8",x"86",x"70",x"4a"),
  1115 => (x"72",x"1e",x"27",x"de"),
  1116 => (x"12",x"00",x"00",x"1e"),
  1117 => (x"27",x"d9",x"00",x"00"),
  1118 => (x"00",x"0f",x"c8",x"86"),
  1119 => (x"72",x"49",x"c1",x"b7"),
  1120 => (x"a9",x"02",x"c0",x"cd"),
  1121 => (x"87",x"27",x"a5",x"10"),
  1122 => (x"00",x"00",x"0f",x"c0"),
  1123 => (x"86",x"c0",x"48",x"c3"),
  1124 => (x"ea",x"87",x"27",x"75"),
  1125 => (x"0e",x"00",x"00",x"0f"),
  1126 => (x"c0",x"86",x"70",x"4c"),
  1127 => (x"74",x"4a",x"cf",x"ff"),
  1128 => (x"ff",x"9a",x"72",x"49"),
  1129 => (x"c6",x"ea",x"b7",x"a9"),
  1130 => (x"02",x"c0",x"dd",x"87"),
  1131 => (x"74",x"1e",x"27",x"87"),
  1132 => (x"12",x"00",x"00",x"1e"),
  1133 => (x"27",x"d9",x"00",x"00"),
  1134 => (x"00",x"0f",x"c8",x"86"),
  1135 => (x"27",x"a5",x"10",x"00"),
  1136 => (x"00",x"0f",x"c0",x"86"),
  1137 => (x"c0",x"48",x"c2",x"f3"),
  1138 => (x"87",x"ff",x"97",x"7b"),
  1139 => (x"c0",x"f1",x"4d",x"27"),
  1140 => (x"c0",x"0f",x"00",x"00"),
  1141 => (x"0f",x"c0",x"86",x"70"),
  1142 => (x"4a",x"72",x"9a",x"02"),
  1143 => (x"c1",x"f7",x"87",x"c0"),
  1144 => (x"1e",x"c0",x"ff",x"f0"),
  1145 => (x"c1",x"fa",x"1e",x"27"),
  1146 => (x"e4",x"0e",x"00",x"00"),
  1147 => (x"0f",x"c8",x"86",x"70"),
  1148 => (x"4c",x"74",x"9c",x"05"),
  1149 => (x"c1",x"cf",x"87",x"74"),
  1150 => (x"1e",x"27",x"9c",x"12"),
  1151 => (x"00",x"00",x"1e",x"27"),
  1152 => (x"d9",x"00",x"00",x"00"),
  1153 => (x"0f",x"c8",x"86",x"ff"),
  1154 => (x"97",x"7b",x"97",x"6b"),
  1155 => (x"48",x"c4",x"a6",x"58"),
  1156 => (x"6e",x"4c",x"c3",x"ff"),
  1157 => (x"9c",x"74",x"1e",x"27"),
  1158 => (x"a8",x"12",x"00",x"00"),
  1159 => (x"1e",x"27",x"d9",x"00"),
  1160 => (x"00",x"00",x"0f",x"c8"),
  1161 => (x"86",x"ff",x"97",x"7b"),
  1162 => (x"ff",x"97",x"7b",x"ff"),
  1163 => (x"97",x"7b",x"ff",x"97"),
  1164 => (x"7b",x"74",x"4a",x"c1"),
  1165 => (x"c0",x"9a",x"72",x"9a"),
  1166 => (x"02",x"c0",x"c5",x"87"),
  1167 => (x"c1",x"48",x"c0",x"fb"),
  1168 => (x"87",x"c0",x"48",x"c0"),
  1169 => (x"f6",x"87",x"74",x"1e"),
  1170 => (x"27",x"b6",x"12",x"00"),
  1171 => (x"00",x"1e",x"27",x"d9"),
  1172 => (x"00",x"00",x"00",x"0f"),
  1173 => (x"c8",x"86",x"75",x"49"),
  1174 => (x"c2",x"b7",x"a9",x"05"),
  1175 => (x"c0",x"d3",x"87",x"27"),
  1176 => (x"c2",x"12",x"00",x"00"),
  1177 => (x"1e",x"27",x"d9",x"00"),
  1178 => (x"00",x"00",x"0f",x"c4"),
  1179 => (x"86",x"c0",x"48",x"c0"),
  1180 => (x"ca",x"87",x"c1",x"8d"),
  1181 => (x"75",x"9d",x"05",x"fd"),
  1182 => (x"d5",x"87",x"c0",x"48"),
  1183 => (x"26",x"26",x"4d",x"26"),
  1184 => (x"4c",x"26",x"4b",x"26"),
  1185 => (x"4a",x"26",x"4f",x"43"),
  1186 => (x"4d",x"44",x"38",x"5f"),
  1187 => (x"34",x"20",x"72",x"65"),
  1188 => (x"73",x"70",x"6f",x"6e"),
  1189 => (x"73",x"65",x"3a",x"20"),
  1190 => (x"25",x"64",x"0a",x"00"),
  1191 => (x"43",x"4d",x"44",x"35"),
  1192 => (x"38",x"20",x"25",x"64"),
  1193 => (x"0a",x"20",x"20",x"00"),
  1194 => (x"43",x"4d",x"44",x"35"),
  1195 => (x"38",x"5f",x"32",x"20"),
  1196 => (x"25",x"64",x"0a",x"20"),
  1197 => (x"20",x"00",x"43",x"4d"),
  1198 => (x"44",x"35",x"38",x"20"),
  1199 => (x"25",x"64",x"0a",x"20"),
  1200 => (x"20",x"00",x"53",x"44"),
  1201 => (x"48",x"43",x"20",x"49"),
  1202 => (x"6e",x"69",x"74",x"69"),
  1203 => (x"61",x"6c",x"69",x"7a"),
  1204 => (x"61",x"74",x"69",x"6f"),
  1205 => (x"6e",x"20",x"65",x"72"),
  1206 => (x"72",x"6f",x"72",x"21"),
  1207 => (x"0a",x"00",x"63",x"6d"),
  1208 => (x"64",x"5f",x"43",x"4d"),
  1209 => (x"44",x"38",x"20",x"72"),
  1210 => (x"65",x"73",x"70",x"6f"),
  1211 => (x"6e",x"73",x"65",x"3a"),
  1212 => (x"20",x"25",x"64",x"0a"),
  1213 => (x"00",x"0e",x"5e",x"5a"),
  1214 => (x"5b",x"5c",x"5d",x"0e"),
  1215 => (x"c0",x"f6",x"e4",x"c0"),
  1216 => (x"c0",x"4d",x"c0",x"f6"),
  1217 => (x"e4",x"c0",x"c4",x"4b"),
  1218 => (x"27",x"e0",x"1a",x"00"),
  1219 => (x"00",x"49",x"c1",x"79"),
  1220 => (x"c0",x"f6",x"e4",x"c0"),
  1221 => (x"c8",x"49",x"c0",x"e0"),
  1222 => (x"51",x"c7",x"4c",x"c3"),
  1223 => (x"97",x"7b",x"27",x"9e"),
  1224 => (x"0f",x"00",x"00",x"0f"),
  1225 => (x"c0",x"86",x"c2",x"97"),
  1226 => (x"7b",x"ff",x"97",x"7d"),
  1227 => (x"c0",x"1e",x"c0",x"e5"),
  1228 => (x"d0",x"c1",x"c0",x"1e"),
  1229 => (x"27",x"e4",x"0e",x"00"),
  1230 => (x"00",x"0f",x"c8",x"86"),
  1231 => (x"70",x"4a",x"72",x"49"),
  1232 => (x"c1",x"b7",x"a9",x"05"),
  1233 => (x"c0",x"c2",x"87",x"c1"),
  1234 => (x"4c",x"74",x"49",x"c2"),
  1235 => (x"b7",x"a9",x"05",x"c0"),
  1236 => (x"c5",x"87",x"c0",x"48"),
  1237 => (x"c0",x"f9",x"87",x"c1"),
  1238 => (x"8c",x"74",x"9c",x"05"),
  1239 => (x"fe",x"fc",x"87",x"27"),
  1240 => (x"43",x"11",x"00",x"00"),
  1241 => (x"0f",x"c0",x"86",x"27"),
  1242 => (x"e0",x"1a",x"00",x"00"),
  1243 => (x"58",x"27",x"e0",x"1a"),
  1244 => (x"00",x"00",x"bf",x"05"),
  1245 => (x"c0",x"d0",x"87",x"c1"),
  1246 => (x"1e",x"c0",x"ff",x"f0"),
  1247 => (x"c1",x"d0",x"1e",x"27"),
  1248 => (x"e4",x"0e",x"00",x"00"),
  1249 => (x"0f",x"c8",x"86",x"ff"),
  1250 => (x"97",x"7d",x"c3",x"53"),
  1251 => (x"ff",x"55",x"c1",x"48"),
  1252 => (x"26",x"4d",x"26",x"4c"),
  1253 => (x"26",x"4b",x"26",x"4a"),
  1254 => (x"26",x"4f",x"1e",x"c0"),
  1255 => (x"48",x"26",x"4f",x"0e"),
  1256 => (x"5e",x"5a",x"5b",x"5c"),
  1257 => (x"5d",x"0e",x"c8",x"8e"),
  1258 => (x"c0",x"e0",x"66",x"4d"),
  1259 => (x"c0",x"f6",x"e4",x"c0"),
  1260 => (x"c0",x"4b",x"76",x"49"),
  1261 => (x"c0",x"79",x"75",x"1e"),
  1262 => (x"c0",x"e0",x"66",x"1e"),
  1263 => (x"27",x"8f",x"14",x"00"),
  1264 => (x"00",x"1e",x"27",x"d9"),
  1265 => (x"00",x"00",x"00",x"0f"),
  1266 => (x"cc",x"86",x"ff",x"97"),
  1267 => (x"7b",x"c0",x"f6",x"e4"),
  1268 => (x"c0",x"c4",x"49",x"c2"),
  1269 => (x"51",x"c0",x"f6",x"e4"),
  1270 => (x"c0",x"c8",x"49",x"c1"),
  1271 => (x"51",x"ff",x"97",x"7b"),
  1272 => (x"dc",x"66",x"1e",x"c0"),
  1273 => (x"ff",x"f0",x"c1",x"d1"),
  1274 => (x"1e",x"27",x"e4",x"0e"),
  1275 => (x"00",x"00",x"0f",x"c8"),
  1276 => (x"86",x"c8",x"a6",x"58"),
  1277 => (x"c4",x"66",x"02",x"c0"),
  1278 => (x"d8",x"87",x"c4",x"66"),
  1279 => (x"1e",x"c0",x"e0",x"66"),
  1280 => (x"1e",x"27",x"6f",x"14"),
  1281 => (x"00",x"00",x"1e",x"27"),
  1282 => (x"d9",x"00",x"00",x"00"),
  1283 => (x"0f",x"cc",x"86",x"c1"),
  1284 => (x"cf",x"87",x"c5",x"ee"),
  1285 => (x"cd",x"df",x"4c",x"ff"),
  1286 => (x"97",x"7b",x"97",x"6b"),
  1287 => (x"48",x"c8",x"a6",x"58"),
  1288 => (x"c4",x"66",x"4a",x"c3"),
  1289 => (x"ff",x"9a",x"72",x"49"),
  1290 => (x"c3",x"fe",x"b7",x"a9"),
  1291 => (x"05",x"c0",x"df",x"87"),
  1292 => (x"c0",x"4a",x"27",x"75"),
  1293 => (x"0e",x"00",x"00",x"0f"),
  1294 => (x"c0",x"86",x"58",x"c4"),
  1295 => (x"85",x"c1",x"82",x"72"),
  1296 => (x"49",x"c2",x"c0",x"b7"),
  1297 => (x"a9",x"04",x"ff",x"e9"),
  1298 => (x"87",x"c1",x"4c",x"76"),
  1299 => (x"49",x"c1",x"79",x"c1"),
  1300 => (x"8c",x"74",x"9c",x"05"),
  1301 => (x"ff",x"c0",x"87",x"ff"),
  1302 => (x"53",x"c0",x"f6",x"e4"),
  1303 => (x"c0",x"c4",x"49",x"c3"),
  1304 => (x"51",x"6e",x"48",x"c8"),
  1305 => (x"86",x"26",x"4d",x"26"),
  1306 => (x"4c",x"26",x"4b",x"26"),
  1307 => (x"4a",x"26",x"4f",x"52"),
  1308 => (x"65",x"61",x"64",x"20"),
  1309 => (x"63",x"6f",x"6d",x"6d"),
  1310 => (x"61",x"6e",x"64",x"20"),
  1311 => (x"66",x"61",x"69",x"6c"),
  1312 => (x"65",x"64",x"20",x"61"),
  1313 => (x"74",x"20",x"25",x"64"),
  1314 => (x"20",x"28",x"25",x"64"),
  1315 => (x"29",x"0a",x"00",x"73"),
  1316 => (x"64",x"5f",x"72",x"65"),
  1317 => (x"61",x"64",x"5f",x"73"),
  1318 => (x"65",x"63",x"74",x"6f"),
  1319 => (x"72",x"20",x"25",x"64"),
  1320 => (x"2c",x"20",x"25",x"64"),
  1321 => (x"0a",x"00",x"1e",x"c0"),
  1322 => (x"f6",x"e8",x"c0",x"c0"),
  1323 => (x"49",x"c4",x"66",x"79"),
  1324 => (x"c4",x"66",x"48",x"26"),
  1325 => (x"4f",x"0e",x"5e",x"5a"),
  1326 => (x"5b",x"5c",x"5d",x"0e"),
  1327 => (x"c8",x"8e",x"c4",x"a6"),
  1328 => (x"49",x"c0",x"79",x"dc"),
  1329 => (x"66",x"4b",x"76",x"49"),
  1330 => (x"23",x"79",x"c0",x"4c"),
  1331 => (x"6e",x"4a",x"d8",x"b7"),
  1332 => (x"2a",x"72",x"4d",x"c3"),
  1333 => (x"ff",x"9d",x"6e",x"48"),
  1334 => (x"c8",x"30",x"c4",x"a6"),
  1335 => (x"58",x"75",x"9d",x"02"),
  1336 => (x"c0",x"e3",x"87",x"75"),
  1337 => (x"1e",x"27",x"a6",x"14"),
  1338 => (x"00",x"00",x"0f",x"c4"),
  1339 => (x"86",x"c4",x"66",x"48"),
  1340 => (x"c1",x"80",x"c8",x"a6"),
  1341 => (x"58",x"c1",x"84",x"74"),
  1342 => (x"49",x"c4",x"b7",x"a9"),
  1343 => (x"04",x"ff",x"cc",x"87"),
  1344 => (x"75",x"9d",x"05",x"ff"),
  1345 => (x"c0",x"87",x"c4",x"66"),
  1346 => (x"48",x"c8",x"86",x"26"),
  1347 => (x"4d",x"26",x"4c",x"26"),
  1348 => (x"4b",x"26",x"4a",x"26"),
  1349 => (x"4f",x"0e",x"5e",x"5a"),
  1350 => (x"5b",x"5c",x"5d",x"0e"),
  1351 => (x"c8",x"8e",x"c0",x"e0"),
  1352 => (x"66",x"4c",x"dc",x"66"),
  1353 => (x"4a",x"76",x"49",x"c0"),
  1354 => (x"79",x"74",x"49",x"c0"),
  1355 => (x"b7",x"a9",x"06",x"c1"),
  1356 => (x"ea",x"87",x"12",x"4b"),
  1357 => (x"c8",x"33",x"c1",x"8c"),
  1358 => (x"74",x"49",x"c0",x"b7"),
  1359 => (x"a9",x"06",x"c0",x"c8"),
  1360 => (x"87",x"12",x"48",x"c8"),
  1361 => (x"a6",x"58",x"c0",x"c5"),
  1362 => (x"87",x"c4",x"a6",x"49"),
  1363 => (x"c0",x"79",x"73",x"4b"),
  1364 => (x"c4",x"66",x"b3",x"c8"),
  1365 => (x"33",x"c1",x"8c",x"74"),
  1366 => (x"49",x"c0",x"b7",x"a9"),
  1367 => (x"06",x"c0",x"c5",x"87"),
  1368 => (x"12",x"4d",x"c0",x"c2"),
  1369 => (x"87",x"c0",x"4d",x"73"),
  1370 => (x"4b",x"75",x"b3",x"c8"),
  1371 => (x"33",x"c1",x"8c",x"74"),
  1372 => (x"49",x"c0",x"b7",x"a9"),
  1373 => (x"06",x"c0",x"c8",x"87"),
  1374 => (x"12",x"48",x"c8",x"a6"),
  1375 => (x"58",x"c0",x"c5",x"87"),
  1376 => (x"c4",x"a6",x"49",x"c0"),
  1377 => (x"79",x"73",x"4b",x"c4"),
  1378 => (x"66",x"b3",x"73",x"48"),
  1379 => (x"6e",x"80",x"c4",x"a6"),
  1380 => (x"58",x"c1",x"8c",x"74"),
  1381 => (x"49",x"c0",x"b7",x"a9"),
  1382 => (x"01",x"fe",x"d6",x"87"),
  1383 => (x"6e",x"48",x"c8",x"86"),
  1384 => (x"26",x"4d",x"26",x"4c"),
  1385 => (x"26",x"4b",x"26",x"4a"),
  1386 => (x"26",x"4f",x"43",x"48"),
  1387 => (x"45",x"43",x"4b",x"53"),
  1388 => (x"55",x"4d",x"42",x"49"),
  1389 => (x"4e",x"00",x"4f",x"53"),
  1390 => (x"44",x"38",x"33",x"32"),
  1391 => (x"30",x"31",x"53",x"59"),
  1392 => (x"53",x"00",x"43",x"61"),
  1393 => (x"6e",x"27",x"74",x"20"),
  1394 => (x"6c",x"6f",x"61",x"64"),
  1395 => (x"20",x"66",x"69",x"72"),
  1396 => (x"6d",x"77",x"61",x"72"),
  1397 => (x"65",x"0a",x"00",x"55"),
  1398 => (x"6e",x"61",x"62",x"6c"),
  1399 => (x"65",x"20",x"74",x"6f"),
  1400 => (x"20",x"6c",x"6f",x"63"),
  1401 => (x"61",x"74",x"65",x"20"),
  1402 => (x"70",x"61",x"72",x"74"),
  1403 => (x"69",x"74",x"69",x"6f"),
  1404 => (x"6e",x"0a",x"00",x"55"),
  1405 => (x"6e",x"61",x"62",x"6c"),
  1406 => (x"65",x"20",x"74",x"6f"),
  1407 => (x"20",x"6c",x"6f",x"63"),
  1408 => (x"61",x"74",x"65",x"20"),
  1409 => (x"70",x"61",x"72",x"74"),
  1410 => (x"69",x"74",x"69",x"6f"),
  1411 => (x"6e",x"0a",x"00",x"48"),
  1412 => (x"75",x"6e",x"74",x"69"),
  1413 => (x"6e",x"67",x"20",x"66"),
  1414 => (x"6f",x"72",x"20",x"70"),
  1415 => (x"61",x"72",x"74",x"69"),
  1416 => (x"74",x"69",x"6f",x"6e"),
  1417 => (x"0a",x"00",x"49",x"6e"),
  1418 => (x"69",x"74",x"69",x"61"),
  1419 => (x"6c",x"69",x"7a",x"69"),
  1420 => (x"6e",x"67",x"20",x"53"),
  1421 => (x"44",x"20",x"63",x"61"),
  1422 => (x"72",x"64",x"0a",x"00"),
  1423 => (x"49",x"6e",x"69",x"74"),
  1424 => (x"69",x"61",x"6c",x"69"),
  1425 => (x"7a",x"69",x"6e",x"67"),
  1426 => (x"20",x"53",x"44",x"20"),
  1427 => (x"63",x"61",x"72",x"64"),
  1428 => (x"0a",x"00",x"46",x"61"),
  1429 => (x"69",x"6c",x"65",x"64"),
  1430 => (x"20",x"74",x"6f",x"20"),
  1431 => (x"69",x"6e",x"69",x"74"),
  1432 => (x"69",x"61",x"6c",x"69"),
  1433 => (x"7a",x"65",x"20",x"53"),
  1434 => (x"44",x"20",x"63",x"61"),
  1435 => (x"72",x"64",x"0a",x"00"),
  1436 => (x"52",x"65",x"61",x"64"),
  1437 => (x"20",x"6f",x"66",x"20"),
  1438 => (x"4d",x"42",x"52",x"20"),
  1439 => (x"66",x"61",x"69",x"6c"),
  1440 => (x"65",x"64",x"0a",x"00"),
  1441 => (x"46",x"41",x"54",x"31"),
  1442 => (x"32",x"20",x"6e",x"6f"),
  1443 => (x"74",x"20",x"73",x"75"),
  1444 => (x"70",x"70",x"6f",x"72"),
  1445 => (x"74",x"65",x"64",x"20"),
  1446 => (x"2d",x"20",x"70",x"6c"),
  1447 => (x"65",x"61",x"73",x"65"),
  1448 => (x"20",x"75",x"73",x"65"),
  1449 => (x"20",x"61",x"20",x"46"),
  1450 => (x"41",x"54",x"31",x"36"),
  1451 => (x"20",x"6f",x"72",x"20"),
  1452 => (x"46",x"41",x"54",x"33"),
  1453 => (x"32",x"20",x"63",x"61"),
  1454 => (x"72",x"64",x"00",x"4e"),
  1455 => (x"6f",x"20",x"70",x"61"),
  1456 => (x"72",x"74",x"69",x"74"),
  1457 => (x"69",x"6f",x"6e",x"20"),
  1458 => (x"73",x"69",x"67",x"6e"),
  1459 => (x"61",x"74",x"75",x"72"),
  1460 => (x"65",x"20",x"66",x"6f"),
  1461 => (x"75",x"6e",x"64",x"0a"),
  1462 => (x"00",x"52",x"65",x"61"),
  1463 => (x"64",x"69",x"6e",x"67"),
  1464 => (x"20",x"62",x"6f",x"6f"),
  1465 => (x"74",x"20",x"73",x"65"),
  1466 => (x"63",x"74",x"6f",x"72"),
  1467 => (x"20",x"25",x"64",x"0a"),
  1468 => (x"00",x"52",x"65",x"61"),
  1469 => (x"64",x"20",x"62",x"6f"),
  1470 => (x"6f",x"74",x"20",x"73"),
  1471 => (x"65",x"63",x"74",x"6f"),
  1472 => (x"72",x"20",x"66",x"72"),
  1473 => (x"6f",x"6d",x"20",x"66"),
  1474 => (x"69",x"72",x"73",x"74"),
  1475 => (x"20",x"70",x"61",x"72"),
  1476 => (x"74",x"69",x"74",x"69"),
  1477 => (x"6f",x"6e",x"0a",x"00"),
  1478 => (x"55",x"6e",x"73",x"75"),
  1479 => (x"70",x"70",x"6f",x"72"),
  1480 => (x"74",x"65",x"64",x"20"),
  1481 => (x"70",x"61",x"72",x"74"),
  1482 => (x"69",x"74",x"69",x"6f"),
  1483 => (x"6e",x"20",x"74",x"79"),
  1484 => (x"70",x"65",x"21",x"0d"),
  1485 => (x"00",x"4f",x"6e",x"6c"),
  1486 => (x"79",x"20",x"46",x"41"),
  1487 => (x"54",x"31",x"36",x"20"),
  1488 => (x"61",x"6e",x"64",x"20"),
  1489 => (x"46",x"41",x"54",x"33"),
  1490 => (x"32",x"20",x"61",x"72"),
  1491 => (x"65",x"20",x"73",x"75"),
  1492 => (x"70",x"70",x"6f",x"72"),
  1493 => (x"74",x"65",x"64",x"0a"),
  1494 => (x"00",x"46",x"41",x"54"),
  1495 => (x"33",x"32",x"20",x"20"),
  1496 => (x"20",x"00",x"52",x"65"),
  1497 => (x"61",x"64",x"69",x"6e"),
  1498 => (x"67",x"20",x"4d",x"42"),
  1499 => (x"52",x"0a",x"00",x"4d"),
  1500 => (x"42",x"52",x"20",x"73"),
  1501 => (x"75",x"63",x"63",x"65"),
  1502 => (x"73",x"73",x"66",x"75"),
  1503 => (x"6c",x"6c",x"79",x"20"),
  1504 => (x"72",x"65",x"61",x"64"),
  1505 => (x"0a",x"00",x"46",x"41"),
  1506 => (x"54",x"31",x"36",x"20"),
  1507 => (x"20",x"20",x"00",x"46"),
  1508 => (x"41",x"54",x"33",x"32"),
  1509 => (x"20",x"20",x"20",x"00"),
  1510 => (x"46",x"41",x"54",x"31"),
  1511 => (x"32",x"20",x"20",x"20"),
  1512 => (x"00",x"50",x"61",x"72"),
  1513 => (x"74",x"69",x"74",x"69"),
  1514 => (x"6f",x"6e",x"63",x"6f"),
  1515 => (x"75",x"6e",x"74",x"20"),
  1516 => (x"25",x"64",x"0a",x"00"),
  1517 => (x"48",x"75",x"6e",x"74"),
  1518 => (x"69",x"6e",x"67",x"20"),
  1519 => (x"66",x"6f",x"72",x"20"),
  1520 => (x"66",x"69",x"6c",x"65"),
  1521 => (x"73",x"79",x"73",x"74"),
  1522 => (x"65",x"6d",x"0a",x"00"),
  1523 => (x"46",x"41",x"54",x"33"),
  1524 => (x"32",x"20",x"20",x"20"),
  1525 => (x"00",x"46",x"41",x"54"),
  1526 => (x"31",x"36",x"20",x"20"),
  1527 => (x"20",x"00",x"47",x"6f"),
  1528 => (x"74",x"20",x"72",x"65"),
  1529 => (x"73",x"75",x"6c",x"74"),
  1530 => (x"20",x"25",x"64",x"20"),
  1531 => (x"0a",x"00",x"64",x"20"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
