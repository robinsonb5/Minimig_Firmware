library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity osdload_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end osdload_ROM;

architecture arch of osdload_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"00",
     2 => x"10",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4f",
     9 => x"f8",
    10 => x"0f",
    11 => x"80",
    12 => x"33",
    13 => x"fc",
    14 => x"55",
    15 => x"55",
    16 => x"00",
    17 => x"00",
    18 => x"04",
    19 => x"12",
    20 => x"61",
    21 => x"00",
    22 => x"02",
    23 => x"80",
    24 => x"66",
    25 => x"50",
    26 => x"33",
    27 => x"fc",
    28 => x"00",
    29 => x"40",
    30 => x"00",
    31 => x"00",
    32 => x"04",
    33 => x"18",
    34 => x"61",
    35 => x"00",
    36 => x"04",
    37 => x"1c",
    38 => x"67",
    39 => x"0c",
    40 => x"42",
    41 => x"79",
    42 => x"00",
    43 => x"00",
    44 => x"04",
    45 => x"18",
    46 => x"61",
    47 => x"00",
    48 => x"04",
    49 => x"10",
    50 => x"66",
    51 => x"2e",
    52 => x"61",
    53 => x"00",
    54 => x"05",
    55 => x"56",
    56 => x"43",
    57 => x"fa",
    58 => x"00",
    59 => x"3c",
    60 => x"61",
    61 => x"00",
    62 => x"05",
    63 => x"9a",
    64 => x"67",
    65 => x"20",
    66 => x"41",
    67 => x"fa",
    68 => x"00",
    69 => x"2c",
    70 => x"61",
    71 => x"00",
    72 => x"03",
    73 => x"7e",
    74 => x"30",
    75 => x"7c",
    76 => x"20",
    77 => x"00",
    78 => x"61",
    79 => x"00",
    80 => x"06",
    81 => x"18",
    82 => x"67",
    83 => x"04",
    84 => x"4e",
    85 => x"f8",
    86 => x"20",
    87 => x"00",
    88 => x"31",
    89 => x"fc",
    90 => x"60",
    91 => x"fe",
    92 => x"20",
    93 => x"00",
    94 => x"4e",
    95 => x"f8",
    96 => x"20",
    97 => x"00",
    98 => x"41",
    99 => x"fa",
   100 => x"00",
   101 => x"08",
   102 => x"61",
   103 => x"00",
   104 => x"03",
   105 => x"5e",
   106 => x"60",
   107 => x"fe",
   108 => x"6e",
   109 => x"6f",
   110 => x"74",
   111 => x"20",
   112 => x"66",
   113 => x"6f",
   114 => x"75",
   115 => x"6e",
   116 => x"64",
   117 => x"20",
   118 => x"4f",
   119 => x"53",
   120 => x"44",
   121 => x"36",
   122 => x"38",
   123 => x"4b",
   124 => x"30",
   125 => x"31",
   126 => x"53",
   127 => x"59",
   128 => x"53",
   129 => x"00",
   130 => x"41",
   131 => x"f8",
   132 => x"10",
   133 => x"00",
   134 => x"0c",
   135 => x"79",
   136 => x"aa",
   137 => x"aa",
   138 => x"00",
   139 => x"00",
   140 => x"04",
   141 => x"12",
   142 => x"66",
   143 => x"0a",
   144 => x"b0",
   145 => x"ba",
   146 => x"03",
   147 => x"82",
   148 => x"66",
   149 => x"04",
   150 => x"70",
   151 => x"00",
   152 => x"4e",
   153 => x"75",
   154 => x"33",
   155 => x"fc",
   156 => x"aa",
   157 => x"aa",
   158 => x"00",
   159 => x"00",
   160 => x"04",
   161 => x"12",
   162 => x"23",
   163 => x"c0",
   164 => x"00",
   165 => x"00",
   166 => x"04",
   167 => x"14",
   168 => x"61",
   169 => x"00",
   170 => x"00",
   171 => x"aa",
   172 => x"66",
   173 => x"4e",
   174 => x"32",
   175 => x"3c",
   176 => x"4e",
   177 => x"20",
   178 => x"12",
   179 => x"bc",
   180 => x"00",
   181 => x"ff",
   182 => x"53",
   183 => x"41",
   184 => x"67",
   185 => x"2e",
   186 => x"30",
   187 => x"11",
   188 => x"12",
   189 => x"bc",
   190 => x"00",
   191 => x"ff",
   192 => x"b0",
   193 => x"3c",
   194 => x"00",
   195 => x"fe",
   196 => x"66",
   197 => x"f0",
   198 => x"32",
   199 => x"3c",
   200 => x"01",
   201 => x"ff",
   202 => x"30",
   203 => x"11",
   204 => x"12",
   205 => x"bc",
   206 => x"00",
   207 => x"ff",
   208 => x"10",
   209 => x"c0",
   210 => x"51",
   211 => x"c9",
   212 => x"ff",
   213 => x"f6",
   214 => x"12",
   215 => x"bc",
   216 => x"00",
   217 => x"ff",
   218 => x"33",
   219 => x"7c",
   220 => x"00",
   221 => x"03",
   222 => x"00",
   223 => x"04",
   224 => x"41",
   225 => x"e8",
   226 => x"fe",
   227 => x"00",
   228 => x"70",
   229 => x"00",
   230 => x"4e",
   231 => x"75",
   232 => x"33",
   233 => x"fc",
   234 => x"55",
   235 => x"55",
   236 => x"00",
   237 => x"00",
   238 => x"04",
   239 => x"12",
   240 => x"41",
   241 => x"fa",
   242 => x"01",
   243 => x"86",
   244 => x"61",
   245 => x"00",
   246 => x"02",
   247 => x"d0",
   248 => x"70",
   249 => x"fe",
   250 => x"4e",
   251 => x"75",
   252 => x"33",
   253 => x"fc",
   254 => x"55",
   255 => x"55",
   256 => x"00",
   257 => x"00",
   258 => x"04",
   259 => x"12",
   260 => x"41",
   261 => x"fa",
   262 => x"01",
   263 => x"5a",
   264 => x"61",
   265 => x"00",
   266 => x"02",
   267 => x"bc",
   268 => x"70",
   269 => x"ff",
   270 => x"4e",
   271 => x"75",
   272 => x"22",
   273 => x"3c",
   274 => x"00",
   275 => x"95",
   276 => x"00",
   277 => x"40",
   278 => x"70",
   279 => x"00",
   280 => x"60",
   281 => x"40",
   282 => x"22",
   283 => x"3c",
   284 => x"00",
   285 => x"ff",
   286 => x"00",
   287 => x"41",
   288 => x"70",
   289 => x"00",
   290 => x"60",
   291 => x"36",
   292 => x"22",
   293 => x"3c",
   294 => x"00",
   295 => x"87",
   296 => x"00",
   297 => x"48",
   298 => x"20",
   299 => x"3c",
   300 => x"00",
   301 => x"00",
   302 => x"01",
   303 => x"aa",
   304 => x"60",
   305 => x"28",
   306 => x"22",
   307 => x"3c",
   308 => x"00",
   309 => x"87",
   310 => x"00",
   311 => x"69",
   312 => x"20",
   313 => x"3c",
   314 => x"40",
   315 => x"00",
   316 => x"00",
   317 => x"00",
   318 => x"60",
   319 => x"1a",
   320 => x"22",
   321 => x"3c",
   322 => x"00",
   323 => x"ff",
   324 => x"00",
   325 => x"77",
   326 => x"70",
   327 => x"00",
   328 => x"60",
   329 => x"10",
   330 => x"22",
   331 => x"3c",
   332 => x"00",
   333 => x"ff",
   334 => x"00",
   335 => x"7a",
   336 => x"70",
   337 => x"00",
   338 => x"60",
   339 => x"06",
   340 => x"22",
   341 => x"3c",
   342 => x"00",
   343 => x"ff",
   344 => x"00",
   345 => x"51",
   346 => x"43",
   347 => x"f9",
   348 => x"00",
   349 => x"da",
   350 => x"40",
   351 => x"00",
   352 => x"12",
   353 => x"bc",
   354 => x"00",
   355 => x"ff",
   356 => x"33",
   357 => x"7c",
   358 => x"00",
   359 => x"02",
   360 => x"00",
   361 => x"04",
   362 => x"12",
   363 => x"81",
   364 => x"48",
   365 => x"41",
   366 => x"4a",
   367 => x"79",
   368 => x"00",
   369 => x"00",
   370 => x"04",
   371 => x"10",
   372 => x"67",
   373 => x"10",
   374 => x"e1",
   375 => x"98",
   376 => x"12",
   377 => x"80",
   378 => x"e1",
   379 => x"98",
   380 => x"12",
   381 => x"80",
   382 => x"e1",
   383 => x"98",
   384 => x"12",
   385 => x"80",
   386 => x"e1",
   387 => x"98",
   388 => x"60",
   389 => x"12",
   390 => x"d0",
   391 => x"80",
   392 => x"48",
   393 => x"40",
   394 => x"12",
   395 => x"80",
   396 => x"48",
   397 => x"40",
   398 => x"e1",
   399 => x"58",
   400 => x"12",
   401 => x"80",
   402 => x"e1",
   403 => x"58",
   404 => x"12",
   405 => x"80",
   406 => x"70",
   407 => x"00",
   408 => x"12",
   409 => x"80",
   410 => x"12",
   411 => x"81",
   412 => x"22",
   413 => x"3c",
   414 => x"00",
   415 => x"00",
   416 => x"9c",
   417 => x"40",
   418 => x"53",
   419 => x"81",
   420 => x"67",
   421 => x"0c",
   422 => x"12",
   423 => x"bc",
   424 => x"00",
   425 => x"ff",
   426 => x"30",
   427 => x"11",
   428 => x"b0",
   429 => x"3c",
   430 => x"00",
   431 => x"ff",
   432 => x"67",
   433 => x"f0",
   434 => x"80",
   435 => x"00",
   436 => x"4e",
   437 => x"75",
   438 => x"d2",
   439 => x"01",
   440 => x"b1",
   441 => x"01",
   442 => x"6a",
   443 => x"04",
   444 => x"0a",
   445 => x"01",
   446 => x"00",
   447 => x"09",
   448 => x"b1",
   449 => x"01",
   450 => x"d0",
   451 => x"00",
   452 => x"d2",
   453 => x"01",
   454 => x"b1",
   455 => x"01",
   456 => x"6a",
   457 => x"04",
   458 => x"0a",
   459 => x"01",
   460 => x"00",
   461 => x"09",
   462 => x"b1",
   463 => x"01",
   464 => x"d0",
   465 => x"00",
   466 => x"d2",
   467 => x"01",
   468 => x"b1",
   469 => x"01",
   470 => x"6a",
   471 => x"04",
   472 => x"0a",
   473 => x"01",
   474 => x"00",
   475 => x"09",
   476 => x"b1",
   477 => x"01",
   478 => x"d0",
   479 => x"00",
   480 => x"d2",
   481 => x"01",
   482 => x"b1",
   483 => x"01",
   484 => x"6a",
   485 => x"04",
   486 => x"0a",
   487 => x"01",
   488 => x"00",
   489 => x"09",
   490 => x"b1",
   491 => x"01",
   492 => x"d0",
   493 => x"00",
   494 => x"d2",
   495 => x"01",
   496 => x"b1",
   497 => x"01",
   498 => x"6a",
   499 => x"04",
   500 => x"0a",
   501 => x"01",
   502 => x"00",
   503 => x"09",
   504 => x"b1",
   505 => x"01",
   506 => x"d0",
   507 => x"00",
   508 => x"d2",
   509 => x"01",
   510 => x"b1",
   511 => x"01",
   512 => x"6a",
   513 => x"04",
   514 => x"0a",
   515 => x"01",
   516 => x"00",
   517 => x"09",
   518 => x"b1",
   519 => x"01",
   520 => x"d0",
   521 => x"00",
   522 => x"d2",
   523 => x"01",
   524 => x"b1",
   525 => x"01",
   526 => x"6a",
   527 => x"04",
   528 => x"0a",
   529 => x"01",
   530 => x"00",
   531 => x"09",
   532 => x"b1",
   533 => x"01",
   534 => x"d0",
   535 => x"00",
   536 => x"d2",
   537 => x"01",
   538 => x"b1",
   539 => x"01",
   540 => x"6a",
   541 => x"04",
   542 => x"0a",
   543 => x"01",
   544 => x"00",
   545 => x"09",
   546 => x"b1",
   547 => x"01",
   548 => x"d0",
   549 => x"00",
   550 => x"4e",
   551 => x"75",
   552 => x"53",
   553 => x"74",
   554 => x"61",
   555 => x"72",
   556 => x"74",
   557 => x"20",
   558 => x"49",
   559 => x"6e",
   560 => x"69",
   561 => x"74",
   562 => x"0d",
   563 => x"0a",
   564 => x"00",
   565 => x"49",
   566 => x"6e",
   567 => x"69",
   568 => x"74",
   569 => x"20",
   570 => x"64",
   571 => x"6f",
   572 => x"6e",
   573 => x"65",
   574 => x"0d",
   575 => x"0a",
   576 => x"00",
   577 => x"49",
   578 => x"6e",
   579 => x"69",
   580 => x"74",
   581 => x"20",
   582 => x"66",
   583 => x"61",
   584 => x"69",
   585 => x"6c",
   586 => x"75",
   587 => x"72",
   588 => x"65",
   589 => x"0d",
   590 => x"0a",
   591 => x"00",
   592 => x"52",
   593 => x"65",
   594 => x"73",
   595 => x"65",
   596 => x"74",
   597 => x"20",
   598 => x"66",
   599 => x"61",
   600 => x"69",
   601 => x"6c",
   602 => x"75",
   603 => x"72",
   604 => x"65",
   605 => x"0d",
   606 => x"0a",
   607 => x"00",
   608 => x"43",
   609 => x"6f",
   610 => x"6d",
   611 => x"6d",
   612 => x"61",
   613 => x"6e",
   614 => x"64",
   615 => x"20",
   616 => x"54",
   617 => x"69",
   618 => x"6d",
   619 => x"65",
   620 => x"6f",
   621 => x"75",
   622 => x"74",
   623 => x"5f",
   624 => x"45",
   625 => x"72",
   626 => x"72",
   627 => x"6f",
   628 => x"72",
   629 => x"0d",
   630 => x"0a",
   631 => x"00",
   632 => x"54",
   633 => x"69",
   634 => x"6d",
   635 => x"65",
   636 => x"6f",
   637 => x"75",
   638 => x"74",
   639 => x"5f",
   640 => x"45",
   641 => x"72",
   642 => x"72",
   643 => x"6f",
   644 => x"72",
   645 => x"0d",
   646 => x"0a",
   647 => x"00",
   648 => x"53",
   649 => x"44",
   650 => x"48",
   651 => x"43",
   652 => x"20",
   653 => x"66",
   654 => x"6f",
   655 => x"75",
   656 => x"6e",
   657 => x"64",
   658 => x"20",
   659 => x"0d",
   660 => x"0a",
   661 => x"00",
   662 => x"33",
   663 => x"fc",
   664 => x"ff",
   665 => x"ff",
   666 => x"00",
   667 => x"00",
   668 => x"04",
   669 => x"10",
   670 => x"43",
   671 => x"f9",
   672 => x"00",
   673 => x"da",
   674 => x"40",
   675 => x"00",
   676 => x"33",
   677 => x"7c",
   678 => x"00",
   679 => x"ff",
   680 => x"00",
   681 => x"04",
   682 => x"33",
   683 => x"7c",
   684 => x"00",
   685 => x"20",
   686 => x"00",
   687 => x"08",
   688 => x"32",
   689 => x"3c",
   690 => x"00",
   691 => x"64",
   692 => x"32",
   693 => x"bc",
   694 => x"ff",
   695 => x"ff",
   696 => x"51",
   697 => x"c9",
   698 => x"ff",
   699 => x"fa",
   700 => x"34",
   701 => x"3c",
   702 => x"00",
   703 => x"32",
   704 => x"61",
   705 => x"00",
   706 => x"fe",
   707 => x"4e",
   708 => x"33",
   709 => x"7c",
   710 => x"00",
   711 => x"03",
   712 => x"00",
   713 => x"04",
   714 => x"b0",
   715 => x"3c",
   716 => x"00",
   717 => x"01",
   718 => x"67",
   719 => x"12",
   720 => x"51",
   721 => x"ca",
   722 => x"ff",
   723 => x"ee",
   724 => x"48",
   725 => x"7a",
   726 => x"ff",
   727 => x"7a",
   728 => x"61",
   729 => x"00",
   730 => x"00",
   731 => x"fa",
   732 => x"58",
   733 => x"8f",
   734 => x"70",
   735 => x"ff",
   736 => x"4e",
   737 => x"75",
   738 => x"22",
   739 => x"3c",
   740 => x"00",
   741 => x"00",
   742 => x"20",
   743 => x"00",
   744 => x"12",
   745 => x"bc",
   746 => x"00",
   747 => x"ff",
   748 => x"53",
   749 => x"81",
   750 => x"66",
   751 => x"f8",
   752 => x"61",
   753 => x"00",
   754 => x"fe",
   755 => x"32",
   756 => x"b0",
   757 => x"3c",
   758 => x"00",
   759 => x"01",
   760 => x"66",
   761 => x"7c",
   762 => x"12",
   763 => x"bc",
   764 => x"00",
   765 => x"ff",
   766 => x"12",
   767 => x"bc",
   768 => x"00",
   769 => x"ff",
   770 => x"12",
   771 => x"bc",
   772 => x"00",
   773 => x"ff",
   774 => x"10",
   775 => x"11",
   776 => x"0c",
   777 => x"00",
   778 => x"00",
   779 => x"01",
   780 => x"66",
   781 => x"68",
   782 => x"12",
   783 => x"bc",
   784 => x"00",
   785 => x"ff",
   786 => x"10",
   787 => x"11",
   788 => x"0c",
   789 => x"00",
   790 => x"00",
   791 => x"aa",
   792 => x"66",
   793 => x"5c",
   794 => x"33",
   795 => x"7c",
   796 => x"00",
   797 => x"03",
   798 => x"00",
   799 => x"04",
   800 => x"48",
   801 => x"7a",
   802 => x"ff",
   803 => x"66",
   804 => x"61",
   805 => x"00",
   806 => x"00",
   807 => x"ae",
   808 => x"58",
   809 => x"8f",
   810 => x"34",
   811 => x"3c",
   812 => x"00",
   813 => x"32",
   814 => x"53",
   815 => x"42",
   816 => x"67",
   817 => x"44",
   818 => x"32",
   819 => x"3c",
   820 => x"07",
   821 => x"d0",
   822 => x"12",
   823 => x"bc",
   824 => x"00",
   825 => x"ff",
   826 => x"51",
   827 => x"c9",
   828 => x"ff",
   829 => x"fa",
   830 => x"61",
   831 => x"00",
   832 => x"fe",
   833 => x"00",
   834 => x"b0",
   835 => x"3c",
   836 => x"00",
   837 => x"01",
   838 => x"66",
   839 => x"e6",
   840 => x"61",
   841 => x"00",
   842 => x"fd",
   843 => x"e8",
   844 => x"66",
   845 => x"e0",
   846 => x"61",
   847 => x"00",
   848 => x"fd",
   849 => x"fa",
   850 => x"66",
   851 => x"da",
   852 => x"12",
   853 => x"bc",
   854 => x"00",
   855 => x"ff",
   856 => x"10",
   857 => x"11",
   858 => x"c0",
   859 => x"3c",
   860 => x"00",
   861 => x"40",
   862 => x"66",
   863 => x"08",
   864 => x"33",
   865 => x"fc",
   866 => x"00",
   867 => x"00",
   868 => x"00",
   869 => x"00",
   870 => x"04",
   871 => x"10",
   872 => x"12",
   873 => x"bc",
   874 => x"00",
   875 => x"ff",
   876 => x"12",
   877 => x"bc",
   878 => x"00",
   879 => x"ff",
   880 => x"12",
   881 => x"bc",
   882 => x"00",
   883 => x"ff",
   884 => x"60",
   885 => x"34",
   886 => x"33",
   887 => x"fc",
   888 => x"00",
   889 => x"00",
   890 => x"00",
   891 => x"00",
   892 => x"04",
   893 => x"10",
   894 => x"34",
   895 => x"3c",
   896 => x"00",
   897 => x"0a",
   898 => x"32",
   899 => x"3c",
   900 => x"07",
   901 => x"d0",
   902 => x"12",
   903 => x"bc",
   904 => x"00",
   905 => x"ff",
   906 => x"51",
   907 => x"c9",
   908 => x"ff",
   909 => x"fa",
   910 => x"61",
   911 => x"00",
   912 => x"fd",
   913 => x"8a",
   914 => x"67",
   915 => x"16",
   916 => x"33",
   917 => x"7c",
   918 => x"00",
   919 => x"03",
   920 => x"00",
   921 => x"04",
   922 => x"51",
   923 => x"ca",
   924 => x"ff",
   925 => x"e6",
   926 => x"48",
   927 => x"7a",
   928 => x"fe",
   929 => x"a1",
   930 => x"61",
   931 => x"30",
   932 => x"58",
   933 => x"8f",
   934 => x"70",
   935 => x"ff",
   936 => x"4e",
   937 => x"75",
   938 => x"33",
   939 => x"7c",
   940 => x"00",
   941 => x"01",
   942 => x"00",
   943 => x"08",
   944 => x"33",
   945 => x"7c",
   946 => x"00",
   947 => x"03",
   948 => x"00",
   949 => x"04",
   950 => x"12",
   951 => x"bc",
   952 => x"00",
   953 => x"ff",
   954 => x"48",
   955 => x"7a",
   956 => x"fe",
   957 => x"79",
   958 => x"61",
   959 => x"14",
   960 => x"58",
   961 => x"8f",
   962 => x"70",
   963 => x"00",
   964 => x"4e",
   965 => x"75",
   966 => x"10",
   967 => x"18",
   968 => x"67",
   969 => x"08",
   970 => x"13",
   971 => x"c0",
   972 => x"00",
   973 => x"da",
   974 => x"80",
   975 => x"00",
   976 => x"60",
   977 => x"f4",
   978 => x"4e",
   979 => x"75",
   980 => x"2f",
   981 => x"08",
   982 => x"20",
   983 => x"6f",
   984 => x"00",
   985 => x"08",
   986 => x"4a",
   987 => x"10",
   988 => x"67",
   989 => x"08",
   990 => x"13",
   991 => x"d8",
   992 => x"00",
   993 => x"da",
   994 => x"80",
   995 => x"00",
   996 => x"60",
   997 => x"f4",
   998 => x"20",
   999 => x"5f",
  1000 => x"4e",
  1001 => x"75",
  1002 => x"00",
  1003 => x"00",
  1004 => x"00",
  1005 => x"00",
  1006 => x"00",
  1007 => x"00",
  1008 => x"00",
  1009 => x"00",
  1010 => x"00",
  1011 => x"00",
  1012 => x"00",
  1013 => x"00",
  1014 => x"00",
  1015 => x"00",
  1016 => x"00",
  1017 => x"00",
  1018 => x"00",
  1019 => x"00",
  1020 => x"00",
  1021 => x"00",
  1022 => x"00",
  1023 => x"00",
  1024 => x"00",
  1025 => x"00",
  1026 => x"00",
  1027 => x"00",
  1028 => x"00",
  1029 => x"00",
  1030 => x"00",
  1031 => x"00",
  1032 => x"00",
  1033 => x"00",
  1034 => x"00",
  1035 => x"00",
  1036 => x"00",
  1037 => x"00",
  1038 => x"00",
  1039 => x"00",
  1040 => x"00",
  1041 => x"00",
  1042 => x"00",
  1043 => x"00",
  1044 => x"00",
  1045 => x"00",
  1046 => x"00",
  1047 => x"00",
  1048 => x"00",
  1049 => x"00",
  1050 => x"00",
  1051 => x"00",
  1052 => x"00",
  1053 => x"00",
  1054 => x"00",
  1055 => x"00",
  1056 => x"00",
  1057 => x"00",
  1058 => x"00",
  1059 => x"00",
  1060 => x"00",
  1061 => x"00",
  1062 => x"00",
  1063 => x"00",
  1064 => x"00",
  1065 => x"00",
  1066 => x"00",
  1067 => x"00",
  1068 => x"00",
  1069 => x"00",
  1070 => x"00",
  1071 => x"00",
  1072 => x"00",
  1073 => x"00",
  1074 => x"00",
  1075 => x"00",
  1076 => x"00",
  1077 => x"00",
  1078 => x"00",
  1079 => x"00",
  1080 => x"00",
  1081 => x"00",
  1082 => x"00",
  1083 => x"00",
  1084 => x"00",
  1085 => x"00",
  1086 => x"00",
  1087 => x"00",
  1088 => x"70",
  1089 => x"00",
  1090 => x"23",
  1091 => x"c0",
  1092 => x"00",
  1093 => x"00",
  1094 => x"04",
  1095 => x"30",
  1096 => x"61",
  1097 => x"00",
  1098 => x"fc",
  1099 => x"38",
  1100 => x"66",
  1101 => x"4a",
  1102 => x"0c",
  1103 => x"28",
  1104 => x"00",
  1105 => x"55",
  1106 => x"01",
  1107 => x"fe",
  1108 => x"66",
  1109 => x"42",
  1110 => x"0c",
  1111 => x"28",
  1112 => x"00",
  1113 => x"aa",
  1114 => x"01",
  1115 => x"ff",
  1116 => x"66",
  1117 => x"3a",
  1118 => x"30",
  1119 => x"3a",
  1120 => x"ff",
  1121 => x"b8",
  1122 => x"c0",
  1123 => x"7c",
  1124 => x"00",
  1125 => x"70",
  1126 => x"b0",
  1127 => x"7c",
  1128 => x"00",
  1129 => x"40",
  1130 => x"64",
  1131 => x"30",
  1132 => x"43",
  1133 => x"e8",
  1134 => x"01",
  1135 => x"be",
  1136 => x"d2",
  1137 => x"c0",
  1138 => x"20",
  1139 => x"29",
  1140 => x"00",
  1141 => x"08",
  1142 => x"e0",
  1143 => x"58",
  1144 => x"48",
  1145 => x"40",
  1146 => x"e0",
  1147 => x"58",
  1148 => x"23",
  1149 => x"c0",
  1150 => x"00",
  1151 => x"00",
  1152 => x"04",
  1153 => x"30",
  1154 => x"61",
  1155 => x"00",
  1156 => x"fb",
  1157 => x"fe",
  1158 => x"66",
  1159 => x"10",
  1160 => x"0c",
  1161 => x"28",
  1162 => x"00",
  1163 => x"55",
  1164 => x"01",
  1165 => x"fe",
  1166 => x"66",
  1167 => x"08",
  1168 => x"0c",
  1169 => x"28",
  1170 => x"00",
  1171 => x"aa",
  1172 => x"01",
  1173 => x"ff",
  1174 => x"67",
  1175 => x"04",
  1176 => x"70",
  1177 => x"ff",
  1178 => x"4e",
  1179 => x"75",
  1180 => x"0c",
  1181 => x"a8",
  1182 => x"46",
  1183 => x"41",
  1184 => x"54",
  1185 => x"31",
  1186 => x"00",
  1187 => x"36",
  1188 => x"66",
  1189 => x"24",
  1190 => x"13",
  1191 => x"fc",
  1192 => x"00",
  1193 => x"0c",
  1194 => x"00",
  1195 => x"00",
  1196 => x"04",
  1197 => x"1a",
  1198 => x"0c",
  1199 => x"a8",
  1200 => x"32",
  1201 => x"20",
  1202 => x"20",
  1203 => x"20",
  1204 => x"00",
  1205 => x"3a",
  1206 => x"67",
  1207 => x"36",
  1208 => x"13",
  1209 => x"fc",
  1210 => x"00",
  1211 => x"10",
  1212 => x"00",
  1213 => x"00",
  1214 => x"04",
  1215 => x"1a",
  1216 => x"0c",
  1217 => x"a8",
  1218 => x"36",
  1219 => x"20",
  1220 => x"20",
  1221 => x"20",
  1222 => x"00",
  1223 => x"3a",
  1224 => x"67",
  1225 => x"24",
  1226 => x"13",
  1227 => x"fc",
  1228 => x"00",
  1229 => x"00",
  1230 => x"00",
  1231 => x"00",
  1232 => x"04",
  1233 => x"1a",
  1234 => x"0c",
  1235 => x"a8",
  1236 => x"46",
  1237 => x"41",
  1238 => x"54",
  1239 => x"33",
  1240 => x"00",
  1241 => x"52",
  1242 => x"66",
  1243 => x"bc",
  1244 => x"0c",
  1245 => x"a8",
  1246 => x"32",
  1247 => x"20",
  1248 => x"20",
  1249 => x"20",
  1250 => x"00",
  1251 => x"56",
  1252 => x"66",
  1253 => x"b2",
  1254 => x"13",
  1255 => x"fc",
  1256 => x"00",
  1257 => x"20",
  1258 => x"00",
  1259 => x"00",
  1260 => x"04",
  1261 => x"1a",
  1262 => x"20",
  1263 => x"28",
  1264 => x"00",
  1265 => x"0a",
  1266 => x"c0",
  1267 => x"bc",
  1268 => x"00",
  1269 => x"ff",
  1270 => x"ff",
  1271 => x"00",
  1272 => x"0c",
  1273 => x"80",
  1274 => x"00",
  1275 => x"00",
  1276 => x"02",
  1277 => x"00",
  1278 => x"66",
  1279 => x"98",
  1280 => x"22",
  1281 => x"3a",
  1282 => x"ff",
  1283 => x"2e",
  1284 => x"30",
  1285 => x"28",
  1286 => x"00",
  1287 => x"0e",
  1288 => x"e0",
  1289 => x"58",
  1290 => x"d2",
  1291 => x"80",
  1292 => x"23",
  1293 => x"c1",
  1294 => x"00",
  1295 => x"00",
  1296 => x"04",
  1297 => x"34",
  1298 => x"0c",
  1299 => x"39",
  1300 => x"00",
  1301 => x"20",
  1302 => x"00",
  1303 => x"00",
  1304 => x"04",
  1305 => x"1a",
  1306 => x"66",
  1307 => x"24",
  1308 => x"20",
  1309 => x"28",
  1310 => x"00",
  1311 => x"2c",
  1312 => x"e0",
  1313 => x"58",
  1314 => x"48",
  1315 => x"40",
  1316 => x"e0",
  1317 => x"58",
  1318 => x"23",
  1319 => x"c0",
  1320 => x"00",
  1321 => x"00",
  1322 => x"04",
  1323 => x"1c",
  1324 => x"20",
  1325 => x"28",
  1326 => x"00",
  1327 => x"24",
  1328 => x"e0",
  1329 => x"58",
  1330 => x"48",
  1331 => x"40",
  1332 => x"e0",
  1333 => x"58",
  1334 => x"d2",
  1335 => x"80",
  1336 => x"53",
  1337 => x"28",
  1338 => x"00",
  1339 => x"10",
  1340 => x"66",
  1341 => x"f8",
  1342 => x"60",
  1343 => x"32",
  1344 => x"70",
  1345 => x"00",
  1346 => x"23",
  1347 => x"c0",
  1348 => x"00",
  1349 => x"00",
  1350 => x"04",
  1351 => x"1c",
  1352 => x"30",
  1353 => x"28",
  1354 => x"00",
  1355 => x"16",
  1356 => x"e0",
  1357 => x"58",
  1358 => x"d2",
  1359 => x"80",
  1360 => x"53",
  1361 => x"28",
  1362 => x"00",
  1363 => x"10",
  1364 => x"66",
  1365 => x"f8",
  1366 => x"23",
  1367 => x"c1",
  1368 => x"00",
  1369 => x"00",
  1370 => x"04",
  1371 => x"20",
  1372 => x"20",
  1373 => x"01",
  1374 => x"10",
  1375 => x"28",
  1376 => x"00",
  1377 => x"12",
  1378 => x"e1",
  1379 => x"48",
  1380 => x"10",
  1381 => x"28",
  1382 => x"00",
  1383 => x"11",
  1384 => x"33",
  1385 => x"c0",
  1386 => x"00",
  1387 => x"00",
  1388 => x"04",
  1389 => x"3e",
  1390 => x"e8",
  1391 => x"48",
  1392 => x"d2",
  1393 => x"80",
  1394 => x"70",
  1395 => x"00",
  1396 => x"10",
  1397 => x"28",
  1398 => x"00",
  1399 => x"0d",
  1400 => x"33",
  1401 => x"c0",
  1402 => x"00",
  1403 => x"00",
  1404 => x"04",
  1405 => x"3c",
  1406 => x"92",
  1407 => x"80",
  1408 => x"92",
  1409 => x"80",
  1410 => x"23",
  1411 => x"c1",
  1412 => x"00",
  1413 => x"00",
  1414 => x"04",
  1415 => x"38",
  1416 => x"70",
  1417 => x"00",
  1418 => x"4e",
  1419 => x"75",
  1420 => x"20",
  1421 => x"3a",
  1422 => x"fe",
  1423 => x"8e",
  1424 => x"23",
  1425 => x"c0",
  1426 => x"00",
  1427 => x"00",
  1428 => x"04",
  1429 => x"24",
  1430 => x"66",
  1431 => x"22",
  1432 => x"42",
  1433 => x"b9",
  1434 => x"00",
  1435 => x"00",
  1436 => x"04",
  1437 => x"24",
  1438 => x"30",
  1439 => x"3a",
  1440 => x"fe",
  1441 => x"9e",
  1442 => x"e8",
  1443 => x"48",
  1444 => x"33",
  1445 => x"c0",
  1446 => x"00",
  1447 => x"00",
  1448 => x"04",
  1449 => x"28",
  1450 => x"20",
  1451 => x"3a",
  1452 => x"fe",
  1453 => x"74",
  1454 => x"23",
  1455 => x"c0",
  1456 => x"00",
  1457 => x"00",
  1458 => x"04",
  1459 => x"2a",
  1460 => x"4e",
  1461 => x"75",
  1462 => x"20",
  1463 => x"3a",
  1464 => x"fe",
  1465 => x"6c",
  1466 => x"32",
  1467 => x"3a",
  1468 => x"fe",
  1469 => x"80",
  1470 => x"33",
  1471 => x"c1",
  1472 => x"00",
  1473 => x"00",
  1474 => x"04",
  1475 => x"28",
  1476 => x"e2",
  1477 => x"49",
  1478 => x"65",
  1479 => x"04",
  1480 => x"e3",
  1481 => x"88",
  1482 => x"60",
  1483 => x"f8",
  1484 => x"d0",
  1485 => x"ba",
  1486 => x"fe",
  1487 => x"6a",
  1488 => x"23",
  1489 => x"c0",
  1490 => x"00",
  1491 => x"00",
  1492 => x"04",
  1493 => x"2a",
  1494 => x"4e",
  1495 => x"75",
  1496 => x"48",
  1497 => x"e7",
  1498 => x"20",
  1499 => x"20",
  1500 => x"24",
  1501 => x"49",
  1502 => x"61",
  1503 => x"00",
  1504 => x"fa",
  1505 => x"a2",
  1506 => x"66",
  1507 => x"78",
  1508 => x"74",
  1509 => x"0f",
  1510 => x"4a",
  1511 => x"10",
  1512 => x"67",
  1513 => x"72",
  1514 => x"70",
  1515 => x"0a",
  1516 => x"12",
  1517 => x"32",
  1518 => x"00",
  1519 => x"00",
  1520 => x"b2",
  1521 => x"30",
  1522 => x"00",
  1523 => x"00",
  1524 => x"67",
  1525 => x"0a",
  1526 => x"d2",
  1527 => x"3c",
  1528 => x"00",
  1529 => x"20",
  1530 => x"b2",
  1531 => x"30",
  1532 => x"00",
  1533 => x"00",
  1534 => x"66",
  1535 => x"36",
  1536 => x"51",
  1537 => x"c8",
  1538 => x"ff",
  1539 => x"ea",
  1540 => x"70",
  1541 => x"00",
  1542 => x"10",
  1543 => x"28",
  1544 => x"00",
  1545 => x"0b",
  1546 => x"33",
  1547 => x"c0",
  1548 => x"00",
  1549 => x"00",
  1550 => x"04",
  1551 => x"2e",
  1552 => x"0c",
  1553 => x"39",
  1554 => x"00",
  1555 => x"20",
  1556 => x"00",
  1557 => x"00",
  1558 => x"04",
  1559 => x"1a",
  1560 => x"66",
  1561 => x"08",
  1562 => x"30",
  1563 => x"28",
  1564 => x"00",
  1565 => x"14",
  1566 => x"e0",
  1567 => x"58",
  1568 => x"48",
  1569 => x"40",
  1570 => x"30",
  1571 => x"28",
  1572 => x"00",
  1573 => x"1a",
  1574 => x"e0",
  1575 => x"58",
  1576 => x"23",
  1577 => x"c0",
  1578 => x"00",
  1579 => x"00",
  1580 => x"04",
  1581 => x"24",
  1582 => x"4c",
  1583 => x"df",
  1584 => x"04",
  1585 => x"04",
  1586 => x"70",
  1587 => x"ff",
  1588 => x"4e",
  1589 => x"75",
  1590 => x"41",
  1591 => x"e8",
  1592 => x"00",
  1593 => x"20",
  1594 => x"51",
  1595 => x"ca",
  1596 => x"ff",
  1597 => x"aa",
  1598 => x"20",
  1599 => x"3a",
  1600 => x"fd",
  1601 => x"ea",
  1602 => x"52",
  1603 => x"80",
  1604 => x"23",
  1605 => x"c0",
  1606 => x"00",
  1607 => x"00",
  1608 => x"04",
  1609 => x"2a",
  1610 => x"53",
  1611 => x"79",
  1612 => x"00",
  1613 => x"00",
  1614 => x"04",
  1615 => x"28",
  1616 => x"66",
  1617 => x"8c",
  1618 => x"61",
  1619 => x"46",
  1620 => x"67",
  1621 => x"06",
  1622 => x"61",
  1623 => x"00",
  1624 => x"ff",
  1625 => x"5e",
  1626 => x"60",
  1627 => x"82",
  1628 => x"4c",
  1629 => x"df",
  1630 => x"04",
  1631 => x"04",
  1632 => x"70",
  1633 => x"00",
  1634 => x"4e",
  1635 => x"75",
  1636 => x"20",
  1637 => x"6f",
  1638 => x"00",
  1639 => x"04",
  1640 => x"61",
  1641 => x"00",
  1642 => x"ff",
  1643 => x"4c",
  1644 => x"61",
  1645 => x"00",
  1646 => x"fa",
  1647 => x"3a",
  1648 => x"66",
  1649 => x"24",
  1650 => x"41",
  1651 => x"e8",
  1652 => x"02",
  1653 => x"00",
  1654 => x"20",
  1655 => x"3a",
  1656 => x"fd",
  1657 => x"b2",
  1658 => x"52",
  1659 => x"80",
  1660 => x"23",
  1661 => x"c0",
  1662 => x"00",
  1663 => x"00",
  1664 => x"04",
  1665 => x"2a",
  1666 => x"53",
  1667 => x"79",
  1668 => x"00",
  1669 => x"00",
  1670 => x"04",
  1671 => x"28",
  1672 => x"66",
  1673 => x"e2",
  1674 => x"2f",
  1675 => x"08",
  1676 => x"61",
  1677 => x"0c",
  1678 => x"20",
  1679 => x"5f",
  1680 => x"66",
  1681 => x"d6",
  1682 => x"20",
  1683 => x"08",
  1684 => x"4e",
  1685 => x"75",
  1686 => x"70",
  1687 => x"00",
  1688 => x"4e",
  1689 => x"75",
  1690 => x"0c",
  1691 => x"39",
  1692 => x"00",
  1693 => x"20",
  1694 => x"00",
  1695 => x"00",
  1696 => x"04",
  1697 => x"1a",
  1698 => x"67",
  1699 => x"38",
  1700 => x"0c",
  1701 => x"39",
  1702 => x"00",
  1703 => x"0c",
  1704 => x"00",
  1705 => x"00",
  1706 => x"04",
  1707 => x"1a",
  1708 => x"67",
  1709 => x"6c",
  1710 => x"20",
  1711 => x"3a",
  1712 => x"fd",
  1713 => x"74",
  1714 => x"e0",
  1715 => x"88",
  1716 => x"d0",
  1717 => x"ba",
  1718 => x"fd",
  1719 => x"7e",
  1720 => x"61",
  1721 => x"00",
  1722 => x"f9",
  1723 => x"c8",
  1724 => x"66",
  1725 => x"58",
  1726 => x"10",
  1727 => x"3a",
  1728 => x"fd",
  1729 => x"67",
  1730 => x"d0",
  1731 => x"40",
  1732 => x"30",
  1733 => x"30",
  1734 => x"00",
  1735 => x"00",
  1736 => x"e0",
  1737 => x"58",
  1738 => x"23",
  1739 => x"c0",
  1740 => x"00",
  1741 => x"00",
  1742 => x"04",
  1743 => x"24",
  1744 => x"80",
  1745 => x"bc",
  1746 => x"ff",
  1747 => x"ff",
  1748 => x"00",
  1749 => x"0f",
  1750 => x"b0",
  1751 => x"7c",
  1752 => x"ff",
  1753 => x"ff",
  1754 => x"4e",
  1755 => x"75",
  1756 => x"20",
  1757 => x"3a",
  1758 => x"fd",
  1759 => x"46",
  1760 => x"ee",
  1761 => x"88",
  1762 => x"d0",
  1763 => x"ba",
  1764 => x"fd",
  1765 => x"50",
  1766 => x"61",
  1767 => x"00",
  1768 => x"f9",
  1769 => x"9a",
  1770 => x"66",
  1771 => x"2a",
  1772 => x"10",
  1773 => x"3a",
  1774 => x"fd",
  1775 => x"39",
  1776 => x"c0",
  1777 => x"7c",
  1778 => x"00",
  1779 => x"7f",
  1780 => x"d0",
  1781 => x"40",
  1782 => x"d0",
  1783 => x"40",
  1784 => x"20",
  1785 => x"30",
  1786 => x"00",
  1787 => x"00",
  1788 => x"e0",
  1789 => x"58",
  1790 => x"48",
  1791 => x"40",
  1792 => x"e0",
  1793 => x"58",
  1794 => x"23",
  1795 => x"c0",
  1796 => x"00",
  1797 => x"00",
  1798 => x"04",
  1799 => x"24",
  1800 => x"80",
  1801 => x"bc",
  1802 => x"f0",
  1803 => x"00",
  1804 => x"00",
  1805 => x"07",
  1806 => x"b0",
  1807 => x"bc",
  1808 => x"ff",
  1809 => x"ff",
  1810 => x"ff",
  1811 => x"ff",
  1812 => x"4e",
  1813 => x"75",
  1814 => x"70",
  1815 => x"00",
  1816 => x"4e",
  1817 => x"75",
  1818 => x"2f",
  1819 => x"02",
  1820 => x"20",
  1821 => x"3a",
  1822 => x"fd",
  1823 => x"06",
  1824 => x"22",
  1825 => x"00",
  1826 => x"d0",
  1827 => x"80",
  1828 => x"d0",
  1829 => x"81",
  1830 => x"22",
  1831 => x"00",
  1832 => x"e0",
  1833 => x"88",
  1834 => x"e4",
  1835 => x"88",
  1836 => x"d0",
  1837 => x"ba",
  1838 => x"fd",
  1839 => x"06",
  1840 => x"24",
  1841 => x"00",
  1842 => x"61",
  1843 => x"00",
  1844 => x"f9",
  1845 => x"4e",
  1846 => x"66",
  1847 => x"52",
  1848 => x"20",
  1849 => x"01",
  1850 => x"e2",
  1851 => x"88",
  1852 => x"c0",
  1853 => x"7c",
  1854 => x"01",
  1855 => x"ff",
  1856 => x"b0",
  1857 => x"7c",
  1858 => x"01",
  1859 => x"ff",
  1860 => x"66",
  1861 => x"14",
  1862 => x"10",
  1863 => x"30",
  1864 => x"00",
  1865 => x"00",
  1866 => x"c1",
  1867 => x"42",
  1868 => x"52",
  1869 => x"80",
  1870 => x"61",
  1871 => x"00",
  1872 => x"f9",
  1873 => x"32",
  1874 => x"66",
  1875 => x"36",
  1876 => x"e1",
  1877 => x"4a",
  1878 => x"14",
  1879 => x"10",
  1880 => x"60",
  1881 => x"0a",
  1882 => x"14",
  1883 => x"30",
  1884 => x"00",
  1885 => x"00",
  1886 => x"e1",
  1887 => x"4a",
  1888 => x"14",
  1889 => x"30",
  1890 => x"00",
  1891 => x"01",
  1892 => x"e1",
  1893 => x"5a",
  1894 => x"c2",
  1895 => x"7c",
  1896 => x"00",
  1897 => x"01",
  1898 => x"67",
  1899 => x"02",
  1900 => x"e8",
  1901 => x"4a",
  1902 => x"c4",
  1903 => x"bc",
  1904 => x"00",
  1905 => x"00",
  1906 => x"0f",
  1907 => x"ff",
  1908 => x"23",
  1909 => x"c2",
  1910 => x"00",
  1911 => x"00",
  1912 => x"04",
  1913 => x"24",
  1914 => x"84",
  1915 => x"bc",
  1916 => x"ff",
  1917 => x"ff",
  1918 => x"f0",
  1919 => x"0f",
  1920 => x"20",
  1921 => x"02",
  1922 => x"24",
  1923 => x"1f",
  1924 => x"b0",
  1925 => x"7c",
  1926 => x"ff",
  1927 => x"ff",
  1928 => x"4e",
  1929 => x"75",
  1930 => x"24",
  1931 => x"1f",
  1932 => x"70",
  1933 => x"00",
  1934 => x"4e",
  1935 => x"75",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

