-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity OSDBoot_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end OSDBoot_ROM;

architecture arch of OSDBoot_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ee040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"88080d80",
     5 => x"04848080",
     6 => x"80950471",
     7 => x"fd060872",
     8 => x"83060981",
     9 => x"05820583",
    10 => x"2b2a83ff",
    11 => x"ff065204",
    12 => x"71fc0608",
    13 => x"72830609",
    14 => x"81058305",
    15 => x"1010102a",
    16 => x"81ff0652",
    17 => x"0471fc06",
    18 => x"08848080",
    19 => x"a1ec7383",
    20 => x"06101005",
    21 => x"08067381",
    22 => x"ff067383",
    23 => x"06098105",
    24 => x"83051010",
    25 => x"102b0772",
    26 => x"fc060c51",
    27 => x"51040284",
    28 => x"05848080",
    29 => x"80880c84",
    30 => x"80808095",
    31 => x"0b848080",
    32 => x"91f10400",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"9fe0e05b",
    36 => x"56807670",
    37 => x"84055808",
    38 => x"715e5e57",
    39 => x"7c708405",
    40 => x"5e085880",
    41 => x"5b77982a",
    42 => x"78882b59",
    43 => x"54738938",
    44 => x"765e8480",
    45 => x"8083e204",
    46 => x"7b802e81",
    47 => x"fd38805c",
    48 => x"7380e42e",
    49 => x"a1387380",
    50 => x"e4268e38",
    51 => x"7380e32e",
    52 => x"819a3884",
    53 => x"808082fa",
    54 => x"047380f3",
    55 => x"2e80f538",
    56 => x"84808082",
    57 => x"fa047584",
    58 => x"1771087e",
    59 => x"5c555752",
    60 => x"7280258e",
    61 => x"38ad5184",
    62 => x"8080919e",
    63 => x"2d720981",
    64 => x"05537280",
    65 => x"2ebe3887",
    66 => x"55729c2a",
    67 => x"73842b54",
    68 => x"5271802e",
    69 => x"83388159",
    70 => x"8972258a",
    71 => x"38b71252",
    72 => x"84808082",
    73 => x"a904b012",
    74 => x"5278802e",
    75 => x"89387151",
    76 => x"84808091",
    77 => x"9e2dff15",
    78 => x"55748025",
    79 => x"cc388480",
    80 => x"8082cc04",
    81 => x"b0518480",
    82 => x"80919e2d",
    83 => x"80538480",
    84 => x"80839304",
    85 => x"75841771",
    86 => x"0870545c",
    87 => x"57528480",
    88 => x"8091b22d",
    89 => x"7b538480",
    90 => x"80839304",
    91 => x"75841771",
    92 => x"08565752",
    93 => x"84808083",
    94 => x"ca04a551",
    95 => x"84808091",
    96 => x"9e2d7351",
    97 => x"84808091",
    98 => x"9e2d8217",
    99 => x"57848080",
   100 => x"83d50472",
   101 => x"ff145452",
   102 => x"807225b9",
   103 => x"38797081",
   104 => x"055b8480",
   105 => x"8080b02d",
   106 => x"70525484",
   107 => x"8080919e",
   108 => x"2d811757",
   109 => x"84808083",
   110 => x"930473a5",
   111 => x"2e098106",
   112 => x"8938815c",
   113 => x"84808083",
   114 => x"d5047351",
   115 => x"84808091",
   116 => x"9e2d8117",
   117 => x"57811b5b",
   118 => x"837b25fd",
   119 => x"c83873fd",
   120 => x"bb387d9f",
   121 => x"e0800c02",
   122 => x"bc050d04",
   123 => x"02f4050d",
   124 => x"7470882a",
   125 => x"83fe8006",
   126 => x"7072982a",
   127 => x"0772882b",
   128 => x"87fc8080",
   129 => x"0673982b",
   130 => x"81f00a06",
   131 => x"71730707",
   132 => x"9fe0800c",
   133 => x"56515351",
   134 => x"028c050d",
   135 => x"0402f805",
   136 => x"0d73882b",
   137 => x"83fe8006",
   138 => x"0284058e",
   139 => x"05848080",
   140 => x"80b02d71",
   141 => x"079fe080",
   142 => x"0c510288",
   143 => x"050d0402",
   144 => x"f8050d73",
   145 => x"70902b71",
   146 => x"902a079f",
   147 => x"e0800c52",
   148 => x"0288050d",
   149 => x"0402f805",
   150 => x"0d735170",
   151 => x"802e8c38",
   152 => x"709fe1a0",
   153 => x"0c800b9f",
   154 => x"e1a80c9f",
   155 => x"e1a80852",
   156 => x"7198389f",
   157 => x"e1a00884",
   158 => x"119fe1a0",
   159 => x"0c70089f",
   160 => x"e1a40c51",
   161 => x"84808085",
   162 => x"94049fe1",
   163 => x"a408882b",
   164 => x"9fe1a40c",
   165 => x"81128306",
   166 => x"9fe1a80c",
   167 => x"9fe1a408",
   168 => x"982c9fe0",
   169 => x"800c0288",
   170 => x"050d0402",
   171 => x"e8050d77",
   172 => x"70525684",
   173 => x"808084d5",
   174 => x"2d9fe080",
   175 => x"08528053",
   176 => x"71802e97",
   177 => x"38811353",
   178 => x"80518480",
   179 => x"8084d52d",
   180 => x"9fe08008",
   181 => x"52848080",
   182 => x"85c00482",
   183 => x"13548155",
   184 => x"900b86e9",
   185 => x"808423a0",
   186 => x"810b86e9",
   187 => x"80802386",
   188 => x"e9808022",
   189 => x"52800b86",
   190 => x"e9808023",
   191 => x"86e98080",
   192 => x"2253800b",
   193 => x"86e98080",
   194 => x"2386e980",
   195 => x"80227083",
   196 => x"ffff0673",
   197 => x"882a7081",
   198 => x"06515451",
   199 => x"5371802e",
   200 => x"81a43874",
   201 => x"802e80e0",
   202 => x"38728280",
   203 => x"862e0981",
   204 => x"06819338",
   205 => x"8055fed5",
   206 => x"ca0b86e9",
   207 => x"80802386",
   208 => x"e9808022",
   209 => x"52810b86",
   210 => x"e9808023",
   211 => x"86e98080",
   212 => x"22527486",
   213 => x"e9808023",
   214 => x"86e98080",
   215 => x"22527386",
   216 => x"e9808023",
   217 => x"86e98080",
   218 => x"22527486",
   219 => x"e9808023",
   220 => x"86e98080",
   221 => x"22527486",
   222 => x"e9808023",
   223 => x"86e98080",
   224 => x"22528480",
   225 => x"8087c604",
   226 => x"73812a82",
   227 => x"80800752",
   228 => x"72722e09",
   229 => x"8106af38",
   230 => x"75518480",
   231 => x"8084d52d",
   232 => x"9fe08008",
   233 => x"53ff1454",
   234 => x"73ff2ea7",
   235 => x"387286e9",
   236 => x"80803486",
   237 => x"e9808033",
   238 => x"5272802e",
   239 => x"e8388051",
   240 => x"84808087",
   241 => x"9a04910b",
   242 => x"86e98084",
   243 => x"23848080",
   244 => x"85e00491",
   245 => x"0b86e980",
   246 => x"8423810b",
   247 => x"9fe0800c",
   248 => x"0298050d",
   249 => x"0402f405",
   250 => x"0d86e980",
   251 => x"8052ff72",
   252 => x"34713353",
   253 => x"ff723472",
   254 => x"882b83fe",
   255 => x"80067233",
   256 => x"7081ff06",
   257 => x"515253ff",
   258 => x"72347271",
   259 => x"07882b72",
   260 => x"337081ff",
   261 => x"06515253",
   262 => x"ff723472",
   263 => x"7107882b",
   264 => x"72337081",
   265 => x"ff067207",
   266 => x"9fe0800c",
   267 => x"5253028c",
   268 => x"050d0402",
   269 => x"ec050d76",
   270 => x"78555574",
   271 => x"86e98080",
   272 => x"349fe1ac",
   273 => x"08853873",
   274 => x"892b5473",
   275 => x"982a5372",
   276 => x"86e98080",
   277 => x"3473902a",
   278 => x"537286e9",
   279 => x"80803473",
   280 => x"882a5372",
   281 => x"86e98080",
   282 => x"347386e9",
   283 => x"80803474",
   284 => x"902a5372",
   285 => x"86e98080",
   286 => x"3486e980",
   287 => x"80337081",
   288 => x"ff065153",
   289 => x"82b8bf54",
   290 => x"7281ff2e",
   291 => x"09810699",
   292 => x"38ff0b86",
   293 => x"e9808034",
   294 => x"86e98080",
   295 => x"337081ff",
   296 => x"06ff1656",
   297 => x"515373e0",
   298 => x"38725284",
   299 => x"8080a1fc",
   300 => x"51848080",
   301 => x"81842d72",
   302 => x"9fe0800c",
   303 => x"0294050d",
   304 => x"0402fc05",
   305 => x"0d81c751",
   306 => x"ff0b86e9",
   307 => x"808034ff",
   308 => x"11517080",
   309 => x"25f23802",
   310 => x"84050d04",
   311 => x"02f0050d",
   312 => x"84808089",
   313 => x"c12d819c",
   314 => x"9f538052",
   315 => x"87fc80f7",
   316 => x"51848080",
   317 => x"88b32d9f",
   318 => x"e0800854",
   319 => x"9fe08008",
   320 => x"812e0981",
   321 => x"0680ea38",
   322 => x"9fe08008",
   323 => x"52848080",
   324 => x"a28c5184",
   325 => x"80808184",
   326 => x"2dff0b86",
   327 => x"e9808034",
   328 => x"820a5284",
   329 => x"9c80e951",
   330 => x"84808088",
   331 => x"b32d9fe0",
   332 => x"8008a138",
   333 => x"9fe08008",
   334 => x"52848080",
   335 => x"a2985184",
   336 => x"80808184",
   337 => x"2dff0b86",
   338 => x"e9808034",
   339 => x"73538480",
   340 => x"808b8904",
   341 => x"9fe08008",
   342 => x"52848080",
   343 => x"a2985184",
   344 => x"80808184",
   345 => x"2d848080",
   346 => x"89c12d84",
   347 => x"80808b82",
   348 => x"049fe080",
   349 => x"08528480",
   350 => x"80a28c51",
   351 => x"84808081",
   352 => x"842dff13",
   353 => x"5372fee2",
   354 => x"38729fe0",
   355 => x"800c0290",
   356 => x"050d0402",
   357 => x"f4050dff",
   358 => x"0b86e980",
   359 => x"80348480",
   360 => x"80a2a451",
   361 => x"84808091",
   362 => x"b22d9353",
   363 => x"805287fc",
   364 => x"80c15184",
   365 => x"808088b3",
   366 => x"2d9fe080",
   367 => x"08a1389f",
   368 => x"e0800852",
   369 => x"848080a2",
   370 => x"b0518480",
   371 => x"8081842d",
   372 => x"ff0b86e9",
   373 => x"80803481",
   374 => x"53848080",
   375 => x"8bfd049f",
   376 => x"e0800852",
   377 => x"848080a2",
   378 => x"b0518480",
   379 => x"8081842d",
   380 => x"84808089",
   381 => x"c12dff13",
   382 => x"5372ffb0",
   383 => x"38729fe0",
   384 => x"800c028c",
   385 => x"050d0402",
   386 => x"f0050d84",
   387 => x"808089c1",
   388 => x"2d83aa52",
   389 => x"849c80c8",
   390 => x"51848080",
   391 => x"88b32d9f",
   392 => x"e080089f",
   393 => x"e0800853",
   394 => x"848080a2",
   395 => x"bc525384",
   396 => x"80808184",
   397 => x"2d72812e",
   398 => x"098106a7",
   399 => x"38848080",
   400 => x"87e52d9f",
   401 => x"e0800883",
   402 => x"ffff0653",
   403 => x"7283aa2e",
   404 => x"ba389fe0",
   405 => x"80085284",
   406 => x"8080a2d4",
   407 => x"51848080",
   408 => x"81842d84",
   409 => x"80808b93",
   410 => x"2d848080",
   411 => x"8d830481",
   412 => x"54848080",
   413 => x"8eb90484",
   414 => x"8080a2ec",
   415 => x"51848080",
   416 => x"81842d80",
   417 => x"54848080",
   418 => x"8eb904ff",
   419 => x"0b86e980",
   420 => x"8034b153",
   421 => x"84808089",
   422 => x"dc2d9fe0",
   423 => x"8008802e",
   424 => x"81883880",
   425 => x"5287fc80",
   426 => x"fa518480",
   427 => x"8088b32d",
   428 => x"9fe08008",
   429 => x"80e3389f",
   430 => x"e0800852",
   431 => x"848080a3",
   432 => x"88518480",
   433 => x"8081842d",
   434 => x"ff0b86e9",
   435 => x"80803486",
   436 => x"e9808033",
   437 => x"7081ff06",
   438 => x"70548480",
   439 => x"80a39453",
   440 => x"51538480",
   441 => x"8081842d",
   442 => x"ff0b86e9",
   443 => x"808034ff",
   444 => x"0b86e980",
   445 => x"8034ff0b",
   446 => x"86e98080",
   447 => x"34ff0b86",
   448 => x"e9808034",
   449 => x"72862a70",
   450 => x"81067056",
   451 => x"51537280",
   452 => x"2ea73884",
   453 => x"80808cef",
   454 => x"049fe080",
   455 => x"08528480",
   456 => x"80a38851",
   457 => x"84808081",
   458 => x"842d7282",
   459 => x"2efec838",
   460 => x"ff135372",
   461 => x"fede3872",
   462 => x"54739fe0",
   463 => x"800c0290",
   464 => x"050d0402",
   465 => x"f4050d81",
   466 => x"0b9fe1ac",
   467 => x"0ca00b86",
   468 => x"e9808834",
   469 => x"830b86e9",
   470 => x"80843484",
   471 => x"808089c1",
   472 => x"2d820b86",
   473 => x"e9808434",
   474 => x"87538052",
   475 => x"84d480c0",
   476 => x"51848080",
   477 => x"88b32d9f",
   478 => x"e0800881",
   479 => x"2e973872",
   480 => x"822e0981",
   481 => x"06893880",
   482 => x"53848080",
   483 => x"8fc704ff",
   484 => x"135372d6",
   485 => x"38848080",
   486 => x"8c872d9f",
   487 => x"e080089f",
   488 => x"e1ac0c81",
   489 => x"5287fc80",
   490 => x"d0518480",
   491 => x"8088b32d",
   492 => x"ff0b86e9",
   493 => x"80803483",
   494 => x"0b86e980",
   495 => x"8434ff0b",
   496 => x"86e98080",
   497 => x"34815372",
   498 => x"9fe0800c",
   499 => x"028c050d",
   500 => x"04800b9f",
   501 => x"e0800c04",
   502 => x"02e4050d",
   503 => x"787a5754",
   504 => x"80765474",
   505 => x"53848080",
   506 => x"a3a45257",
   507 => x"84808081",
   508 => x"842dff0b",
   509 => x"86e98080",
   510 => x"34820b86",
   511 => x"e9808434",
   512 => x"810b86e9",
   513 => x"808834ff",
   514 => x"0b86e980",
   515 => x"80347352",
   516 => x"87fc80d1",
   517 => x"51848080",
   518 => x"88b32d80",
   519 => x"dbc6df55",
   520 => x"9fe08008",
   521 => x"772e9a38",
   522 => x"9fe08008",
   523 => x"53735284",
   524 => x"8080a3bc",
   525 => x"51848080",
   526 => x"81842d84",
   527 => x"80809194",
   528 => x"04ff0b86",
   529 => x"e9808034",
   530 => x"86e98080",
   531 => x"337081ff",
   532 => x"06515473",
   533 => x"81fe2e09",
   534 => x"8106a438",
   535 => x"80ff5484",
   536 => x"808087e5",
   537 => x"2d9fe080",
   538 => x"08767084",
   539 => x"05580cff",
   540 => x"14547380",
   541 => x"25e93881",
   542 => x"57848080",
   543 => x"918604ff",
   544 => x"155574ff",
   545 => x"bc38ff0b",
   546 => x"86e98080",
   547 => x"34830b86",
   548 => x"e9808434",
   549 => x"769fe080",
   550 => x"0c029c05",
   551 => x"0d0402fc",
   552 => x"050d7270",
   553 => x"86ea8080",
   554 => x"0c9fe080",
   555 => x"0c028405",
   556 => x"0d0402ec",
   557 => x"050d8077",
   558 => x"56547470",
   559 => x"84055608",
   560 => x"51805370",
   561 => x"982a7188",
   562 => x"2b525271",
   563 => x"802e9838",
   564 => x"7186ea80",
   565 => x"800c8114",
   566 => x"81145454",
   567 => x"837325e3",
   568 => x"38848080",
   569 => x"91ba0473",
   570 => x"9fe0800c",
   571 => x"0294050d",
   572 => x"0402f805",
   573 => x"0d848080",
   574 => x"a3dc5184",
   575 => x"808091b2",
   576 => x"2d848080",
   577 => x"8ec32d9f",
   578 => x"e0800880",
   579 => x"2ebb3884",
   580 => x"8080a3f4",
   581 => x"51848080",
   582 => x"91b22d84",
   583 => x"808093ab",
   584 => x"2d805284",
   585 => x"8080a48c",
   586 => x"51848080",
   587 => x"9fa22d9f",
   588 => x"e0800880",
   589 => x"2e873884",
   590 => x"8080808c",
   591 => x"2d848080",
   592 => x"a4985184",
   593 => x"808091b2",
   594 => x"2d848080",
   595 => x"a4b05184",
   596 => x"808091b2",
   597 => x"2d800b9f",
   598 => x"e0800c02",
   599 => x"88050d04",
   600 => x"02e8050d",
   601 => x"77797b58",
   602 => x"55558053",
   603 => x"727625af",
   604 => x"38747081",
   605 => x"05568480",
   606 => x"8080b02d",
   607 => x"74708105",
   608 => x"56848080",
   609 => x"80b02d52",
   610 => x"5271712e",
   611 => x"89388151",
   612 => x"84808093",
   613 => x"a1048113",
   614 => x"53848080",
   615 => x"92ec0480",
   616 => x"51709fe0",
   617 => x"800c0298",
   618 => x"050d0402",
   619 => x"d8050dff",
   620 => x"0b9fe5d8",
   621 => x"0c800b9f",
   622 => x"e5ec0c84",
   623 => x"8080a4d0",
   624 => x"51848080",
   625 => x"91b22d9f",
   626 => x"e1c45280",
   627 => x"51848080",
   628 => x"8fd82d9f",
   629 => x"e0800854",
   630 => x"9fe08008",
   631 => x"95388480",
   632 => x"80a4e051",
   633 => x"84808091",
   634 => x"b22d7355",
   635 => x"8480809b",
   636 => x"86048480",
   637 => x"80a4f451",
   638 => x"84808091",
   639 => x"b22d8056",
   640 => x"810b9fe1",
   641 => x"b80c8853",
   642 => x"848080a5",
   643 => x"8c529fe1",
   644 => x"fa518480",
   645 => x"8092e02d",
   646 => x"9fe08008",
   647 => x"762e0981",
   648 => x"0689389f",
   649 => x"e080089f",
   650 => x"e1b80c88",
   651 => x"53848080",
   652 => x"a598529f",
   653 => x"e2965184",
   654 => x"808092e0",
   655 => x"2d9fe080",
   656 => x"0889389f",
   657 => x"e080089f",
   658 => x"e1b80c9f",
   659 => x"e1b80852",
   660 => x"848080a5",
   661 => x"a4518480",
   662 => x"8081842d",
   663 => x"9fe1b808",
   664 => x"802e81c1",
   665 => x"389fe58a",
   666 => x"0b848080",
   667 => x"80b02d9f",
   668 => x"e58b0b84",
   669 => x"808080b0",
   670 => x"2d71982b",
   671 => x"71902b07",
   672 => x"9fe58c0b",
   673 => x"84808080",
   674 => x"b02d7088",
   675 => x"2b72079f",
   676 => x"e58d0b84",
   677 => x"808080b0",
   678 => x"2d71079f",
   679 => x"e5c20b84",
   680 => x"808080b0",
   681 => x"2d9fe5c3",
   682 => x"0b848080",
   683 => x"80b02d71",
   684 => x"882b0753",
   685 => x"5f54525a",
   686 => x"56575573",
   687 => x"81abaa2e",
   688 => x"09810694",
   689 => x"38755184",
   690 => x"808083ec",
   691 => x"2d9fe080",
   692 => x"08568480",
   693 => x"8095f104",
   694 => x"7382d4d5",
   695 => x"2e933884",
   696 => x"8080a5b8",
   697 => x"51848080",
   698 => x"91b22d84",
   699 => x"808097f0",
   700 => x"04755284",
   701 => x"8080a5d8",
   702 => x"51848080",
   703 => x"81842d9f",
   704 => x"e1c45275",
   705 => x"51848080",
   706 => x"8fd82d9f",
   707 => x"e0800855",
   708 => x"9fe08008",
   709 => x"802e84ee",
   710 => x"38848080",
   711 => x"a5f05184",
   712 => x"808091b2",
   713 => x"2d848080",
   714 => x"a6985184",
   715 => x"80808184",
   716 => x"2d885384",
   717 => x"8080a598",
   718 => x"529fe296",
   719 => x"51848080",
   720 => x"92e02d9f",
   721 => x"e080088d",
   722 => x"38810b9f",
   723 => x"e5ec0c84",
   724 => x"80809781",
   725 => x"04885384",
   726 => x"8080a58c",
   727 => x"529fe1fa",
   728 => x"51848080",
   729 => x"92e02d9f",
   730 => x"e0800880",
   731 => x"2e933884",
   732 => x"8080a6b0",
   733 => x"51848080",
   734 => x"81842d84",
   735 => x"808097f0",
   736 => x"049fe5c2",
   737 => x"0b848080",
   738 => x"80b02d54",
   739 => x"7380d52e",
   740 => x"09810680",
   741 => x"db389fe5",
   742 => x"c30b8480",
   743 => x"8080b02d",
   744 => x"547381aa",
   745 => x"2e098106",
   746 => x"80c63880",
   747 => x"0b9fe1c4",
   748 => x"0b848080",
   749 => x"80b02d56",
   750 => x"547481e9",
   751 => x"2e833881",
   752 => x"547481eb",
   753 => x"2e8c3880",
   754 => x"5573752e",
   755 => x"09810683",
   756 => x"b5389fe1",
   757 => x"cf0b8480",
   758 => x"8080b02d",
   759 => x"55749138",
   760 => x"9fe1d00b",
   761 => x"84808080",
   762 => x"b02d5473",
   763 => x"822e8938",
   764 => x"80558480",
   765 => x"809b8604",
   766 => x"9fe1d10b",
   767 => x"84808080",
   768 => x"b02d709f",
   769 => x"e5f40cff",
   770 => x"059fe5e8",
   771 => x"0c9fe1d2",
   772 => x"0b848080",
   773 => x"80b02d9f",
   774 => x"e1d30b84",
   775 => x"808080b0",
   776 => x"2d587605",
   777 => x"77828029",
   778 => x"05709fe5",
   779 => x"dc0c9fe1",
   780 => x"d40b8480",
   781 => x"8080b02d",
   782 => x"709fe5d4",
   783 => x"0c9fe5ec",
   784 => x"08595758",
   785 => x"76802e81",
   786 => x"d7388853",
   787 => x"848080a5",
   788 => x"98529fe2",
   789 => x"96518480",
   790 => x"8092e02d",
   791 => x"9fe08008",
   792 => x"82a4389f",
   793 => x"e5f40870",
   794 => x"842b9fe5",
   795 => x"c40c709f",
   796 => x"e5f00c9f",
   797 => x"e1e90b84",
   798 => x"808080b0",
   799 => x"2d9fe1e8",
   800 => x"0b848080",
   801 => x"80b02d71",
   802 => x"82802905",
   803 => x"9fe1ea0b",
   804 => x"84808080",
   805 => x"b02d7084",
   806 => x"80802912",
   807 => x"9fe1eb0b",
   808 => x"84808080",
   809 => x"b02d7081",
   810 => x"800a2912",
   811 => x"709fe1bc",
   812 => x"0c9fe5d4",
   813 => x"0871299f",
   814 => x"e5dc0805",
   815 => x"709fe5fc",
   816 => x"0c9fe1f1",
   817 => x"0b848080",
   818 => x"80b02d9f",
   819 => x"e1f00b84",
   820 => x"808080b0",
   821 => x"2d718280",
   822 => x"29059fe1",
   823 => x"f20b8480",
   824 => x"8080b02d",
   825 => x"70848080",
   826 => x"29129fe1",
   827 => x"f30b8480",
   828 => x"8080b02d",
   829 => x"70982b81",
   830 => x"f00a0672",
   831 => x"05709fe1",
   832 => x"c00cfe11",
   833 => x"7e297705",
   834 => x"9fe5e40c",
   835 => x"52595243",
   836 => x"545e5152",
   837 => x"59525d57",
   838 => x"59578480",
   839 => x"809b8404",
   840 => x"9fe1d60b",
   841 => x"84808080",
   842 => x"b02d9fe1",
   843 => x"d50b8480",
   844 => x"8080b02d",
   845 => x"71828029",
   846 => x"05709fe5",
   847 => x"c40c70a0",
   848 => x"2983ff05",
   849 => x"70892a70",
   850 => x"9fe5f00c",
   851 => x"9fe1db0b",
   852 => x"84808080",
   853 => x"b02d9fe1",
   854 => x"da0b8480",
   855 => x"8080b02d",
   856 => x"71828029",
   857 => x"05709fe1",
   858 => x"bc0c7b71",
   859 => x"291e709f",
   860 => x"e5e40c7d",
   861 => x"9fe1c00c",
   862 => x"73059fe5",
   863 => x"fc0c555e",
   864 => x"51515555",
   865 => x"8155749f",
   866 => x"e0800c02",
   867 => x"a8050d04",
   868 => x"02ec050d",
   869 => x"7670872c",
   870 => x"7180ff06",
   871 => x"5755539f",
   872 => x"e5ec088a",
   873 => x"3872882c",
   874 => x"7381ff06",
   875 => x"5654739f",
   876 => x"e5d8082e",
   877 => x"a4389fe1",
   878 => x"c4529fe5",
   879 => x"dc081451",
   880 => x"8480808f",
   881 => x"d82d9fe0",
   882 => x"8008539f",
   883 => x"e0800880",
   884 => x"2e80c938",
   885 => x"739fe5d8",
   886 => x"0c9fe5ec",
   887 => x"08802ea0",
   888 => x"38748429",
   889 => x"9fe1c405",
   890 => x"70085253",
   891 => x"84808083",
   892 => x"ec2d9fe0",
   893 => x"8008f00a",
   894 => x"06558480",
   895 => x"809c9a04",
   896 => x"74109fe1",
   897 => x"c4057084",
   898 => x"8080809b",
   899 => x"2d525384",
   900 => x"8080849d",
   901 => x"2d9fe080",
   902 => x"08557453",
   903 => x"729fe080",
   904 => x"0c029405",
   905 => x"0d0402cc",
   906 => x"050d7e60",
   907 => x"5e5b8056",
   908 => x"ff0b9fe5",
   909 => x"d80c9fe1",
   910 => x"c0089fe5",
   911 => x"e4085657",
   912 => x"9fe5ec08",
   913 => x"762e8e38",
   914 => x"9fe5f408",
   915 => x"842b5984",
   916 => x"80809cdc",
   917 => x"049fe5f0",
   918 => x"08842b59",
   919 => x"805a7979",
   920 => x"2781e838",
   921 => x"798f06a0",
   922 => x"17575473",
   923 => x"a2387452",
   924 => x"848080a6",
   925 => x"d0518480",
   926 => x"8081842d",
   927 => x"9fe1c452",
   928 => x"74518115",
   929 => x"55848080",
   930 => x"8fd82d9f",
   931 => x"e1c45680",
   932 => x"76848080",
   933 => x"80b02d55",
   934 => x"5873782e",
   935 => x"83388158",
   936 => x"7381e52e",
   937 => x"819c3881",
   938 => x"70790655",
   939 => x"5c73802e",
   940 => x"8190388b",
   941 => x"16848080",
   942 => x"80b02d98",
   943 => x"06587781",
   944 => x"81388b53",
   945 => x"7c527551",
   946 => x"84808092",
   947 => x"e02d9fe0",
   948 => x"800880ee",
   949 => x"389c1608",
   950 => x"51848080",
   951 => x"83ec2d9f",
   952 => x"e0800884",
   953 => x"1c0c9a16",
   954 => x"84808080",
   955 => x"9b2d5184",
   956 => x"8080849d",
   957 => x"2d9fe080",
   958 => x"089fe080",
   959 => x"0855559f",
   960 => x"e5ec0880",
   961 => x"2e9f3894",
   962 => x"16848080",
   963 => x"809b2d51",
   964 => x"84808084",
   965 => x"9d2d9fe0",
   966 => x"8008902b",
   967 => x"83fff00a",
   968 => x"06701651",
   969 => x"5473881c",
   970 => x"0c777b0c",
   971 => x"7c528480",
   972 => x"80a6f051",
   973 => x"84808081",
   974 => x"842d7b54",
   975 => x"8480809f",
   976 => x"9804811a",
   977 => x"5a848080",
   978 => x"9cde049f",
   979 => x"e5ec0880",
   980 => x"2e80c338",
   981 => x"76518480",
   982 => x"809b902d",
   983 => x"9fe08008",
   984 => x"9fe08008",
   985 => x"53848080",
   986 => x"a7845257",
   987 => x"84808081",
   988 => x"842d7680",
   989 => x"fffffff8",
   990 => x"06547380",
   991 => x"fffffff8",
   992 => x"2e9438fe",
   993 => x"179fe5f4",
   994 => x"08299fe5",
   995 => x"fc080555",
   996 => x"8480809c",
   997 => x"dc048054",
   998 => x"739fe080",
   999 => x"0c02b405",
  1000 => x"0d0402e4",
  1001 => x"050d787a",
  1002 => x"71549fe5",
  1003 => x"c8535555",
  1004 => x"8480809c",
  1005 => x"a62d9fe0",
  1006 => x"800881ff",
  1007 => x"06537280",
  1008 => x"2e80fe38",
  1009 => x"848080a7",
  1010 => x"9c518480",
  1011 => x"8091b22d",
  1012 => x"9fe5cc08",
  1013 => x"83ff0589",
  1014 => x"2a578070",
  1015 => x"56567577",
  1016 => x"2580fd38",
  1017 => x"9fe5d008",
  1018 => x"fe059fe5",
  1019 => x"f408299f",
  1020 => x"e5fc0811",
  1021 => x"769fe5e8",
  1022 => x"08060575",
  1023 => x"54525384",
  1024 => x"80808fd8",
  1025 => x"2d9fe080",
  1026 => x"08802e80",
  1027 => x"c8388115",
  1028 => x"709fe5e8",
  1029 => x"08065455",
  1030 => x"7294389f",
  1031 => x"e5d00851",
  1032 => x"8480809b",
  1033 => x"902d9fe0",
  1034 => x"80089fe5",
  1035 => x"d00c8480",
  1036 => x"14811757",
  1037 => x"54767624",
  1038 => x"ffaa3884",
  1039 => x"8080a0e0",
  1040 => x"04745284",
  1041 => x"8080a7b8",
  1042 => x"51848080",
  1043 => x"81842d84",
  1044 => x"8080a0e2",
  1045 => x"049fe080",
  1046 => x"08538480",
  1047 => x"80a0e204",
  1048 => x"8153729f",
  1049 => x"e0800c02",
  1050 => x"9c050d04",
  1051 => x"9fe08c08",
  1052 => x"029fe08c",
  1053 => x"0cff3d0d",
  1054 => x"800b9fe0",
  1055 => x"8c08fc05",
  1056 => x"0c9fe08c",
  1057 => x"08880508",
  1058 => x"8106ff11",
  1059 => x"7009709f",
  1060 => x"e08c088c",
  1061 => x"0508069f",
  1062 => x"e08c08fc",
  1063 => x"0508119f",
  1064 => x"e08c08fc",
  1065 => x"050c9fe0",
  1066 => x"8c088805",
  1067 => x"08812a9f",
  1068 => x"e08c0888",
  1069 => x"050c9fe0",
  1070 => x"8c088c05",
  1071 => x"08109fe0",
  1072 => x"8c088c05",
  1073 => x"0c515151",
  1074 => x"519fe08c",
  1075 => x"08880508",
  1076 => x"802e8438",
  1077 => x"ffab399f",
  1078 => x"e08c08fc",
  1079 => x"0508709f",
  1080 => x"e0800c51",
  1081 => x"833d0d9f",
  1082 => x"e08c0c04",
  1083 => x"00ffffff",
  1084 => x"ff00ffff",
  1085 => x"ffff00ff",
  1086 => x"ffffff00",
  1087 => x"476f7420",
  1088 => x"72657375",
  1089 => x"6c742025",
  1090 => x"64200a00",
  1091 => x"434d4435",
  1092 => x"35202564",
  1093 => x"0a000000",
  1094 => x"434d4434",
  1095 => x"31202564",
  1096 => x"0a000000",
  1097 => x"436d645f",
  1098 => x"696e6974",
  1099 => x"0a000000",
  1100 => x"696e6974",
  1101 => x"2025640a",
  1102 => x"20200000",
  1103 => x"636d645f",
  1104 => x"434d4438",
  1105 => x"20726573",
  1106 => x"706f6e73",
  1107 => x"653a2025",
  1108 => x"640a0000",
  1109 => x"434d4438",
  1110 => x"5f342072",
  1111 => x"6573706f",
  1112 => x"6e73653a",
  1113 => x"2025640a",
  1114 => x"00000000",
  1115 => x"53444843",
  1116 => x"20496e69",
  1117 => x"7469616c",
  1118 => x"697a6174",
  1119 => x"696f6e20",
  1120 => x"6572726f",
  1121 => x"72210a00",
  1122 => x"434d4435",
  1123 => x"38202564",
  1124 => x"0a202000",
  1125 => x"434d4435",
  1126 => x"385f3220",
  1127 => x"25640a20",
  1128 => x"20000000",
  1129 => x"73645f72",
  1130 => x"6561645f",
  1131 => x"73656374",
  1132 => x"6f722025",
  1133 => x"642c2025",
  1134 => x"640a0000",
  1135 => x"52656164",
  1136 => x"20636f6d",
  1137 => x"6d616e64",
  1138 => x"20666169",
  1139 => x"6c656420",
  1140 => x"61742025",
  1141 => x"64202825",
  1142 => x"64290a00",
  1143 => x"496e6974",
  1144 => x"69616c69",
  1145 => x"7a696e67",
  1146 => x"20534420",
  1147 => x"63617264",
  1148 => x"0a000000",
  1149 => x"48756e74",
  1150 => x"696e6720",
  1151 => x"666f7220",
  1152 => x"70617274",
  1153 => x"6974696f",
  1154 => x"6e0a0000",
  1155 => x"4f53445a",
  1156 => x"50553031",
  1157 => x"53595300",
  1158 => x"43616e27",
  1159 => x"74206c6f",
  1160 => x"61642066",
  1161 => x"69726d77",
  1162 => x"6172650a",
  1163 => x"00000000",
  1164 => x"4661696c",
  1165 => x"65642074",
  1166 => x"6f20696e",
  1167 => x"69746961",
  1168 => x"6c697a65",
  1169 => x"20534420",
  1170 => x"63617264",
  1171 => x"0a000000",
  1172 => x"52656164",
  1173 => x"696e6720",
  1174 => x"4d42520a",
  1175 => x"00000000",
  1176 => x"52656164",
  1177 => x"206f6620",
  1178 => x"4d425220",
  1179 => x"6661696c",
  1180 => x"65640a00",
  1181 => x"4d425220",
  1182 => x"73756363",
  1183 => x"65737366",
  1184 => x"756c6c79",
  1185 => x"20726561",
  1186 => x"640a0000",
  1187 => x"46415431",
  1188 => x"36202020",
  1189 => x"00000000",
  1190 => x"46415433",
  1191 => x"32202020",
  1192 => x"00000000",
  1193 => x"50617274",
  1194 => x"6974696f",
  1195 => x"6e636f75",
  1196 => x"6e742025",
  1197 => x"640a0000",
  1198 => x"4e6f2070",
  1199 => x"61727469",
  1200 => x"74696f6e",
  1201 => x"20736967",
  1202 => x"6e617475",
  1203 => x"72652066",
  1204 => x"6f756e64",
  1205 => x"0a000000",
  1206 => x"52656164",
  1207 => x"696e6720",
  1208 => x"626f6f74",
  1209 => x"20736563",
  1210 => x"746f7220",
  1211 => x"25640a00",
  1212 => x"52656164",
  1213 => x"20626f6f",
  1214 => x"74207365",
  1215 => x"63746f72",
  1216 => x"2066726f",
  1217 => x"6d206669",
  1218 => x"72737420",
  1219 => x"70617274",
  1220 => x"6974696f",
  1221 => x"6e0a0000",
  1222 => x"48756e74",
  1223 => x"696e6720",
  1224 => x"666f7220",
  1225 => x"66696c65",
  1226 => x"73797374",
  1227 => x"656d0a00",
  1228 => x"556e7375",
  1229 => x"70706f72",
  1230 => x"74656420",
  1231 => x"70617274",
  1232 => x"6974696f",
  1233 => x"6e207479",
  1234 => x"7065210d",
  1235 => x"00000000",
  1236 => x"52656164",
  1237 => x"696e6720",
  1238 => x"64697265",
  1239 => x"63746f72",
  1240 => x"79207365",
  1241 => x"63746f72",
  1242 => x"2025640a",
  1243 => x"00000000",
  1244 => x"66696c65",
  1245 => x"20222573",
  1246 => x"2220666f",
  1247 => x"756e640d",
  1248 => x"00000000",
  1249 => x"47657446",
  1250 => x"41544c69",
  1251 => x"6e6b2072",
  1252 => x"65747572",
  1253 => x"6e656420",
  1254 => x"25640a00",
  1255 => x"4f70656e",
  1256 => x"65642066",
  1257 => x"696c652c",
  1258 => x"206c6f61",
  1259 => x"64696e67",
  1260 => x"2e2e2e0a",
  1261 => x"00000000",
  1262 => x"43616e27",
  1263 => x"74206f70",
  1264 => x"656e2025",
  1265 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

