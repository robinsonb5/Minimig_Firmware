-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity OSDBoot_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end OSDBoot_ROM;

architecture arch of OSDBoot_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"0b0b9fe0",
     9 => x"80080b0b",
    10 => x"9fe08408",
    11 => x"0b0b9fe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b0b9f",
    15 => x"e0880c0b",
    16 => x"0b9fe084",
    17 => x"0c0b0b9f",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080a1ec",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"9fe08070",
    57 => x"9fe68027",
    58 => x"8e388071",
    59 => x"70840553",
    60 => x"0c848080",
    61 => x"81e30484",
    62 => x"8080808c",
    63 => x"51848080",
    64 => x"92f00402",
    65 => x"c4050d02",
    66 => x"80c0059f",
    67 => x"e0e05b56",
    68 => x"80767084",
    69 => x"05580871",
    70 => x"5e5e577c",
    71 => x"7084055e",
    72 => x"0858805b",
    73 => x"77982a78",
    74 => x"882b5954",
    75 => x"73893876",
    76 => x"5e848080",
    77 => x"84e1047b",
    78 => x"802e81fd",
    79 => x"38805c73",
    80 => x"80e42ea1",
    81 => x"387380e4",
    82 => x"268e3873",
    83 => x"80e32e81",
    84 => x"9a388480",
    85 => x"8083f904",
    86 => x"7380f32e",
    87 => x"80f53884",
    88 => x"808083f9",
    89 => x"04758417",
    90 => x"71087e5c",
    91 => x"55575272",
    92 => x"80258e38",
    93 => x"ad518480",
    94 => x"80929d2d",
    95 => x"72098105",
    96 => x"5372802e",
    97 => x"be388755",
    98 => x"729c2a73",
    99 => x"842b5452",
   100 => x"71802e83",
   101 => x"38815989",
   102 => x"72258a38",
   103 => x"b7125284",
   104 => x"808083a8",
   105 => x"04b01252",
   106 => x"78802e89",
   107 => x"38715184",
   108 => x"8080929d",
   109 => x"2dff1555",
   110 => x"748025cc",
   111 => x"38848080",
   112 => x"83cb04b0",
   113 => x"51848080",
   114 => x"929d2d80",
   115 => x"53848080",
   116 => x"84920475",
   117 => x"84177108",
   118 => x"70545c57",
   119 => x"52848080",
   120 => x"92b12d7b",
   121 => x"53848080",
   122 => x"84920475",
   123 => x"84177108",
   124 => x"56575284",
   125 => x"808084c9",
   126 => x"04a55184",
   127 => x"8080929d",
   128 => x"2d735184",
   129 => x"8080929d",
   130 => x"2d821757",
   131 => x"84808084",
   132 => x"d40472ff",
   133 => x"14545280",
   134 => x"7225b938",
   135 => x"79708105",
   136 => x"5b848080",
   137 => x"80f52d70",
   138 => x"52548480",
   139 => x"80929d2d",
   140 => x"81175784",
   141 => x"80808492",
   142 => x"0473a52e",
   143 => x"09810689",
   144 => x"38815c84",
   145 => x"808084d4",
   146 => x"04735184",
   147 => x"8080929d",
   148 => x"2d811757",
   149 => x"811b5b83",
   150 => x"7b25fdc8",
   151 => x"3873fdbb",
   152 => x"387d9fe0",
   153 => x"800c02bc",
   154 => x"050d0402",
   155 => x"f4050d74",
   156 => x"70882a83",
   157 => x"fe800670",
   158 => x"72982a07",
   159 => x"72882b87",
   160 => x"fc808006",
   161 => x"73982b81",
   162 => x"f00a0671",
   163 => x"7307079f",
   164 => x"e0800c56",
   165 => x"51535102",
   166 => x"8c050d04",
   167 => x"02f8050d",
   168 => x"73882b83",
   169 => x"fe800602",
   170 => x"84058e05",
   171 => x"84808080",
   172 => x"f52d7107",
   173 => x"9fe0800c",
   174 => x"51028805",
   175 => x"0d0402f8",
   176 => x"050d7370",
   177 => x"902b7190",
   178 => x"2a079fe0",
   179 => x"800c5202",
   180 => x"88050d04",
   181 => x"02f8050d",
   182 => x"73517080",
   183 => x"2e8c3870",
   184 => x"9fe1a00c",
   185 => x"800b9fe1",
   186 => x"a80c9fe1",
   187 => x"a8085271",
   188 => x"98389fe1",
   189 => x"a0088411",
   190 => x"9fe1a00c",
   191 => x"70089fe1",
   192 => x"a40c5184",
   193 => x"80808693",
   194 => x"049fe1a4",
   195 => x"08882b9f",
   196 => x"e1a40c81",
   197 => x"1283069f",
   198 => x"e1a80c9f",
   199 => x"e1a40898",
   200 => x"2c9fe080",
   201 => x"0c028805",
   202 => x"0d0402e8",
   203 => x"050d7770",
   204 => x"52568480",
   205 => x"8085d42d",
   206 => x"9fe08008",
   207 => x"52805371",
   208 => x"802e9738",
   209 => x"81135380",
   210 => x"51848080",
   211 => x"85d42d9f",
   212 => x"e0800852",
   213 => x"84808086",
   214 => x"bf048213",
   215 => x"54815590",
   216 => x"0b86e980",
   217 => x"8423a081",
   218 => x"0b86e980",
   219 => x"802386e9",
   220 => x"80802252",
   221 => x"800b86e9",
   222 => x"80802386",
   223 => x"e9808022",
   224 => x"53800b86",
   225 => x"e9808023",
   226 => x"86e98080",
   227 => x"227083ff",
   228 => x"ff067388",
   229 => x"2a708106",
   230 => x"51545153",
   231 => x"71802e81",
   232 => x"a4387480",
   233 => x"2e80e038",
   234 => x"72828086",
   235 => x"2e098106",
   236 => x"81933880",
   237 => x"55fed5ca",
   238 => x"0b86e980",
   239 => x"802386e9",
   240 => x"80802252",
   241 => x"810b86e9",
   242 => x"80802386",
   243 => x"e9808022",
   244 => x"527486e9",
   245 => x"80802386",
   246 => x"e9808022",
   247 => x"527386e9",
   248 => x"80802386",
   249 => x"e9808022",
   250 => x"527486e9",
   251 => x"80802386",
   252 => x"e9808022",
   253 => x"527486e9",
   254 => x"80802386",
   255 => x"e9808022",
   256 => x"52848080",
   257 => x"88c50473",
   258 => x"812a8280",
   259 => x"80075272",
   260 => x"722e0981",
   261 => x"06af3875",
   262 => x"51848080",
   263 => x"85d42d9f",
   264 => x"e0800853",
   265 => x"ff145473",
   266 => x"ff2ea738",
   267 => x"7286e980",
   268 => x"803486e9",
   269 => x"80803352",
   270 => x"72802ee8",
   271 => x"38805184",
   272 => x"80808899",
   273 => x"04910b86",
   274 => x"e9808423",
   275 => x"84808086",
   276 => x"df04910b",
   277 => x"86e98084",
   278 => x"23810b9f",
   279 => x"e0800c02",
   280 => x"98050d04",
   281 => x"02f4050d",
   282 => x"86e98080",
   283 => x"52ff7234",
   284 => x"713353ff",
   285 => x"72347288",
   286 => x"2b83fe80",
   287 => x"06723370",
   288 => x"81ff0651",
   289 => x"5253ff72",
   290 => x"34727107",
   291 => x"882b7233",
   292 => x"7081ff06",
   293 => x"515253ff",
   294 => x"72347271",
   295 => x"07882b72",
   296 => x"337081ff",
   297 => x"0672079f",
   298 => x"e0800c52",
   299 => x"53028c05",
   300 => x"0d0402ec",
   301 => x"050d7678",
   302 => x"55557486",
   303 => x"e9808034",
   304 => x"9fe1ac08",
   305 => x"85387389",
   306 => x"2b547398",
   307 => x"2a537286",
   308 => x"e9808034",
   309 => x"73902a53",
   310 => x"7286e980",
   311 => x"80347388",
   312 => x"2a537286",
   313 => x"e9808034",
   314 => x"7386e980",
   315 => x"80347490",
   316 => x"2a537286",
   317 => x"e9808034",
   318 => x"86e98080",
   319 => x"337081ff",
   320 => x"06515382",
   321 => x"b8bf5472",
   322 => x"81ff2e09",
   323 => x"81069938",
   324 => x"ff0b86e9",
   325 => x"80803486",
   326 => x"e9808033",
   327 => x"7081ff06",
   328 => x"ff165651",
   329 => x"5373e038",
   330 => x"72528480",
   331 => x"80a1fc51",
   332 => x"84808082",
   333 => x"832d729f",
   334 => x"e0800c02",
   335 => x"94050d04",
   336 => x"02fc050d",
   337 => x"81c751ff",
   338 => x"0b86e980",
   339 => x"8034ff11",
   340 => x"51708025",
   341 => x"f2380284",
   342 => x"050d0402",
   343 => x"f0050d84",
   344 => x"80808ac0",
   345 => x"2d819c9f",
   346 => x"53805287",
   347 => x"fc80f751",
   348 => x"84808089",
   349 => x"b22d9fe0",
   350 => x"8008549f",
   351 => x"e0800881",
   352 => x"2e098106",
   353 => x"80ea389f",
   354 => x"e0800852",
   355 => x"848080a2",
   356 => x"8c518480",
   357 => x"8082832d",
   358 => x"ff0b86e9",
   359 => x"80803482",
   360 => x"0a52849c",
   361 => x"80e95184",
   362 => x"808089b2",
   363 => x"2d9fe080",
   364 => x"08a1389f",
   365 => x"e0800852",
   366 => x"848080a2",
   367 => x"98518480",
   368 => x"8082832d",
   369 => x"ff0b86e9",
   370 => x"80803473",
   371 => x"53848080",
   372 => x"8c88049f",
   373 => x"e0800852",
   374 => x"848080a2",
   375 => x"98518480",
   376 => x"8082832d",
   377 => x"8480808a",
   378 => x"c02d8480",
   379 => x"808c8104",
   380 => x"9fe08008",
   381 => x"52848080",
   382 => x"a28c5184",
   383 => x"80808283",
   384 => x"2dff1353",
   385 => x"72fee238",
   386 => x"729fe080",
   387 => x"0c029005",
   388 => x"0d0402f4",
   389 => x"050dff0b",
   390 => x"86e98080",
   391 => x"34848080",
   392 => x"a2a45184",
   393 => x"808092b1",
   394 => x"2d935380",
   395 => x"5287fc80",
   396 => x"c1518480",
   397 => x"8089b22d",
   398 => x"9fe08008",
   399 => x"a1389fe0",
   400 => x"80085284",
   401 => x"8080a2b0",
   402 => x"51848080",
   403 => x"82832dff",
   404 => x"0b86e980",
   405 => x"80348153",
   406 => x"8480808c",
   407 => x"fc049fe0",
   408 => x"80085284",
   409 => x"8080a2b0",
   410 => x"51848080",
   411 => x"82832d84",
   412 => x"80808ac0",
   413 => x"2dff1353",
   414 => x"72ffb038",
   415 => x"729fe080",
   416 => x"0c028c05",
   417 => x"0d0402f0",
   418 => x"050d8480",
   419 => x"808ac02d",
   420 => x"83aa5284",
   421 => x"9c80c851",
   422 => x"84808089",
   423 => x"b22d9fe0",
   424 => x"80089fe0",
   425 => x"80085384",
   426 => x"8080a2bc",
   427 => x"52538480",
   428 => x"8082832d",
   429 => x"72812e09",
   430 => x"8106a738",
   431 => x"84808088",
   432 => x"e42d9fe0",
   433 => x"800883ff",
   434 => x"ff065372",
   435 => x"83aa2eba",
   436 => x"389fe080",
   437 => x"08528480",
   438 => x"80a2d451",
   439 => x"84808082",
   440 => x"832d8480",
   441 => x"808c922d",
   442 => x"8480808e",
   443 => x"82048154",
   444 => x"8480808f",
   445 => x"b8048480",
   446 => x"80a2ec51",
   447 => x"84808082",
   448 => x"832d8054",
   449 => x"8480808f",
   450 => x"b804ff0b",
   451 => x"86e98080",
   452 => x"34b15384",
   453 => x"80808adb",
   454 => x"2d9fe080",
   455 => x"08802e81",
   456 => x"88388052",
   457 => x"87fc80fa",
   458 => x"51848080",
   459 => x"89b22d9f",
   460 => x"e0800880",
   461 => x"e3389fe0",
   462 => x"80085284",
   463 => x"8080a388",
   464 => x"51848080",
   465 => x"82832dff",
   466 => x"0b86e980",
   467 => x"803486e9",
   468 => x"80803370",
   469 => x"81ff0670",
   470 => x"54848080",
   471 => x"a3945351",
   472 => x"53848080",
   473 => x"82832dff",
   474 => x"0b86e980",
   475 => x"8034ff0b",
   476 => x"86e98080",
   477 => x"34ff0b86",
   478 => x"e9808034",
   479 => x"ff0b86e9",
   480 => x"80803472",
   481 => x"862a7081",
   482 => x"06705651",
   483 => x"5372802e",
   484 => x"a7388480",
   485 => x"808dee04",
   486 => x"9fe08008",
   487 => x"52848080",
   488 => x"a3885184",
   489 => x"80808283",
   490 => x"2d72822e",
   491 => x"fec838ff",
   492 => x"135372fe",
   493 => x"de387254",
   494 => x"739fe080",
   495 => x"0c029005",
   496 => x"0d0402f4",
   497 => x"050d810b",
   498 => x"9fe1ac0c",
   499 => x"a00b86e9",
   500 => x"80883483",
   501 => x"0b86e980",
   502 => x"84348480",
   503 => x"808ac02d",
   504 => x"820b86e9",
   505 => x"80843487",
   506 => x"53805284",
   507 => x"d480c051",
   508 => x"84808089",
   509 => x"b22d9fe0",
   510 => x"8008812e",
   511 => x"97387282",
   512 => x"2e098106",
   513 => x"89388053",
   514 => x"84808090",
   515 => x"c604ff13",
   516 => x"5372d638",
   517 => x"8480808d",
   518 => x"862d9fe0",
   519 => x"80089fe1",
   520 => x"ac0c8152",
   521 => x"87fc80d0",
   522 => x"51848080",
   523 => x"89b22dff",
   524 => x"0b86e980",
   525 => x"8034830b",
   526 => x"86e98084",
   527 => x"34ff0b86",
   528 => x"e9808034",
   529 => x"8153729f",
   530 => x"e0800c02",
   531 => x"8c050d04",
   532 => x"800b9fe0",
   533 => x"800c0402",
   534 => x"e4050d78",
   535 => x"7a575480",
   536 => x"76547453",
   537 => x"848080a3",
   538 => x"a4525784",
   539 => x"80808283",
   540 => x"2dff0b86",
   541 => x"e9808034",
   542 => x"820b86e9",
   543 => x"80843481",
   544 => x"0b86e980",
   545 => x"8834ff0b",
   546 => x"86e98080",
   547 => x"34735287",
   548 => x"fc80d151",
   549 => x"84808089",
   550 => x"b22d80db",
   551 => x"c6df559f",
   552 => x"e0800877",
   553 => x"2e9a389f",
   554 => x"e0800853",
   555 => x"73528480",
   556 => x"80a3bc51",
   557 => x"84808082",
   558 => x"832d8480",
   559 => x"80929304",
   560 => x"ff0b86e9",
   561 => x"80803486",
   562 => x"e9808033",
   563 => x"7081ff06",
   564 => x"51547381",
   565 => x"fe2e0981",
   566 => x"06a43880",
   567 => x"ff548480",
   568 => x"8088e42d",
   569 => x"9fe08008",
   570 => x"76708405",
   571 => x"580cff14",
   572 => x"54738025",
   573 => x"e9388157",
   574 => x"84808092",
   575 => x"8504ff15",
   576 => x"5574ffbc",
   577 => x"38ff0b86",
   578 => x"e9808034",
   579 => x"830b86e9",
   580 => x"80843476",
   581 => x"9fe0800c",
   582 => x"029c050d",
   583 => x"0402fc05",
   584 => x"0d727086",
   585 => x"ea80800c",
   586 => x"9fe0800c",
   587 => x"0284050d",
   588 => x"0402ec05",
   589 => x"0d807756",
   590 => x"54747084",
   591 => x"05560851",
   592 => x"80537098",
   593 => x"2a71882b",
   594 => x"52527180",
   595 => x"2e983871",
   596 => x"86ea8080",
   597 => x"0c811481",
   598 => x"14545483",
   599 => x"7325e338",
   600 => x"84808092",
   601 => x"b904739f",
   602 => x"e0800c02",
   603 => x"94050d04",
   604 => x"02f8050d",
   605 => x"848080a3",
   606 => x"dc518480",
   607 => x"8092b12d",
   608 => x"8480808f",
   609 => x"c22d9fe0",
   610 => x"8008802e",
   611 => x"bb388480",
   612 => x"80a3f451",
   613 => x"84808092",
   614 => x"b12d8480",
   615 => x"8094aa2d",
   616 => x"80528480",
   617 => x"80a48c51",
   618 => x"848080a0",
   619 => x"a12d9fe0",
   620 => x"8008802e",
   621 => x"87388480",
   622 => x"8080932d",
   623 => x"848080a4",
   624 => x"98518480",
   625 => x"8092b12d",
   626 => x"848080a4",
   627 => x"b0518480",
   628 => x"8092b12d",
   629 => x"800b9fe0",
   630 => x"800c0288",
   631 => x"050d0402",
   632 => x"e8050d77",
   633 => x"797b5855",
   634 => x"55805372",
   635 => x"7625af38",
   636 => x"74708105",
   637 => x"56848080",
   638 => x"80f52d74",
   639 => x"70810556",
   640 => x"84808080",
   641 => x"f52d5252",
   642 => x"71712e89",
   643 => x"38815184",
   644 => x"808094a0",
   645 => x"04811353",
   646 => x"84808093",
   647 => x"eb048051",
   648 => x"709fe080",
   649 => x"0c029805",
   650 => x"0d0402d8",
   651 => x"050dff0b",
   652 => x"9fe5d80c",
   653 => x"800b9fe5",
   654 => x"ec0c8480",
   655 => x"80a4d051",
   656 => x"84808092",
   657 => x"b12d9fe1",
   658 => x"c4528051",
   659 => x"84808090",
   660 => x"d72d9fe0",
   661 => x"8008549f",
   662 => x"e0800895",
   663 => x"38848080",
   664 => x"a4e05184",
   665 => x"808092b1",
   666 => x"2d735584",
   667 => x"80809c85",
   668 => x"04848080",
   669 => x"a4f45184",
   670 => x"808092b1",
   671 => x"2d805681",
   672 => x"0b9fe1b8",
   673 => x"0c885384",
   674 => x"8080a58c",
   675 => x"529fe1fa",
   676 => x"51848080",
   677 => x"93df2d9f",
   678 => x"e0800876",
   679 => x"2e098106",
   680 => x"89389fe0",
   681 => x"80089fe1",
   682 => x"b80c8853",
   683 => x"848080a5",
   684 => x"98529fe2",
   685 => x"96518480",
   686 => x"8093df2d",
   687 => x"9fe08008",
   688 => x"89389fe0",
   689 => x"80089fe1",
   690 => x"b80c9fe1",
   691 => x"b8085284",
   692 => x"8080a5a4",
   693 => x"51848080",
   694 => x"82832d9f",
   695 => x"e1b80880",
   696 => x"2e81c138",
   697 => x"9fe58a0b",
   698 => x"84808080",
   699 => x"f52d9fe5",
   700 => x"8b0b8480",
   701 => x"8080f52d",
   702 => x"71982b71",
   703 => x"902b079f",
   704 => x"e58c0b84",
   705 => x"808080f5",
   706 => x"2d70882b",
   707 => x"72079fe5",
   708 => x"8d0b8480",
   709 => x"8080f52d",
   710 => x"71079fe5",
   711 => x"c20b8480",
   712 => x"8080f52d",
   713 => x"9fe5c30b",
   714 => x"84808080",
   715 => x"f52d7188",
   716 => x"2b07535f",
   717 => x"54525a56",
   718 => x"57557381",
   719 => x"abaa2e09",
   720 => x"81069438",
   721 => x"75518480",
   722 => x"8084eb2d",
   723 => x"9fe08008",
   724 => x"56848080",
   725 => x"96f00473",
   726 => x"82d4d52e",
   727 => x"93388480",
   728 => x"80a5b851",
   729 => x"84808092",
   730 => x"b12d8480",
   731 => x"8098ef04",
   732 => x"75528480",
   733 => x"80a5d851",
   734 => x"84808082",
   735 => x"832d9fe1",
   736 => x"c4527551",
   737 => x"84808090",
   738 => x"d72d9fe0",
   739 => x"8008559f",
   740 => x"e0800880",
   741 => x"2e84ee38",
   742 => x"848080a5",
   743 => x"f0518480",
   744 => x"8092b12d",
   745 => x"848080a6",
   746 => x"98518480",
   747 => x"8082832d",
   748 => x"88538480",
   749 => x"80a59852",
   750 => x"9fe29651",
   751 => x"84808093",
   752 => x"df2d9fe0",
   753 => x"80088d38",
   754 => x"810b9fe5",
   755 => x"ec0c8480",
   756 => x"80988004",
   757 => x"88538480",
   758 => x"80a58c52",
   759 => x"9fe1fa51",
   760 => x"84808093",
   761 => x"df2d9fe0",
   762 => x"8008802e",
   763 => x"93388480",
   764 => x"80a6b051",
   765 => x"84808082",
   766 => x"832d8480",
   767 => x"8098ef04",
   768 => x"9fe5c20b",
   769 => x"84808080",
   770 => x"f52d5473",
   771 => x"80d52e09",
   772 => x"810680db",
   773 => x"389fe5c3",
   774 => x"0b848080",
   775 => x"80f52d54",
   776 => x"7381aa2e",
   777 => x"09810680",
   778 => x"c638800b",
   779 => x"9fe1c40b",
   780 => x"84808080",
   781 => x"f52d5654",
   782 => x"7481e92e",
   783 => x"83388154",
   784 => x"7481eb2e",
   785 => x"8c388055",
   786 => x"73752e09",
   787 => x"810683b5",
   788 => x"389fe1cf",
   789 => x"0b848080",
   790 => x"80f52d55",
   791 => x"7491389f",
   792 => x"e1d00b84",
   793 => x"808080f5",
   794 => x"2d547382",
   795 => x"2e893880",
   796 => x"55848080",
   797 => x"9c85049f",
   798 => x"e1d10b84",
   799 => x"808080f5",
   800 => x"2d709fe5",
   801 => x"f40cff05",
   802 => x"9fe5e80c",
   803 => x"9fe1d20b",
   804 => x"84808080",
   805 => x"f52d9fe1",
   806 => x"d30b8480",
   807 => x"8080f52d",
   808 => x"58760577",
   809 => x"82802905",
   810 => x"709fe5dc",
   811 => x"0c9fe1d4",
   812 => x"0b848080",
   813 => x"80f52d70",
   814 => x"9fe5d40c",
   815 => x"9fe5ec08",
   816 => x"59575876",
   817 => x"802e81d7",
   818 => x"38885384",
   819 => x"8080a598",
   820 => x"529fe296",
   821 => x"51848080",
   822 => x"93df2d9f",
   823 => x"e0800882",
   824 => x"a4389fe5",
   825 => x"f4087084",
   826 => x"2b9fe5c4",
   827 => x"0c709fe5",
   828 => x"f00c9fe1",
   829 => x"e90b8480",
   830 => x"8080f52d",
   831 => x"9fe1e80b",
   832 => x"84808080",
   833 => x"f52d7182",
   834 => x"8029059f",
   835 => x"e1ea0b84",
   836 => x"808080f5",
   837 => x"2d708480",
   838 => x"8029129f",
   839 => x"e1eb0b84",
   840 => x"808080f5",
   841 => x"2d708180",
   842 => x"0a291270",
   843 => x"9fe1bc0c",
   844 => x"9fe5d408",
   845 => x"71299fe5",
   846 => x"dc080570",
   847 => x"9fe5fc0c",
   848 => x"9fe1f10b",
   849 => x"84808080",
   850 => x"f52d9fe1",
   851 => x"f00b8480",
   852 => x"8080f52d",
   853 => x"71828029",
   854 => x"059fe1f2",
   855 => x"0b848080",
   856 => x"80f52d70",
   857 => x"84808029",
   858 => x"129fe1f3",
   859 => x"0b848080",
   860 => x"80f52d70",
   861 => x"982b81f0",
   862 => x"0a067205",
   863 => x"709fe1c0",
   864 => x"0cfe117e",
   865 => x"2977059f",
   866 => x"e5e40c52",
   867 => x"59524354",
   868 => x"5e515259",
   869 => x"525d5759",
   870 => x"57848080",
   871 => x"9c83049f",
   872 => x"e1d60b84",
   873 => x"808080f5",
   874 => x"2d9fe1d5",
   875 => x"0b848080",
   876 => x"80f52d71",
   877 => x"82802905",
   878 => x"709fe5c4",
   879 => x"0c70a029",
   880 => x"83ff0570",
   881 => x"892a709f",
   882 => x"e5f00c9f",
   883 => x"e1db0b84",
   884 => x"808080f5",
   885 => x"2d9fe1da",
   886 => x"0b848080",
   887 => x"80f52d71",
   888 => x"82802905",
   889 => x"709fe1bc",
   890 => x"0c7b7129",
   891 => x"1e709fe5",
   892 => x"e40c7d9f",
   893 => x"e1c00c73",
   894 => x"059fe5fc",
   895 => x"0c555e51",
   896 => x"51555581",
   897 => x"55749fe0",
   898 => x"800c02a8",
   899 => x"050d0402",
   900 => x"ec050d76",
   901 => x"70872c71",
   902 => x"80ff0657",
   903 => x"55539fe5",
   904 => x"ec088a38",
   905 => x"72882c73",
   906 => x"81ff0656",
   907 => x"54739fe5",
   908 => x"d8082ea4",
   909 => x"389fe1c4",
   910 => x"529fe5dc",
   911 => x"08145184",
   912 => x"808090d7",
   913 => x"2d9fe080",
   914 => x"08539fe0",
   915 => x"8008802e",
   916 => x"80c93873",
   917 => x"9fe5d80c",
   918 => x"9fe5ec08",
   919 => x"802ea038",
   920 => x"7484299f",
   921 => x"e1c40570",
   922 => x"08525384",
   923 => x"808084eb",
   924 => x"2d9fe080",
   925 => x"08f00a06",
   926 => x"55848080",
   927 => x"9d990474",
   928 => x"109fe1c4",
   929 => x"05708480",
   930 => x"8080e02d",
   931 => x"52538480",
   932 => x"80859c2d",
   933 => x"9fe08008",
   934 => x"55745372",
   935 => x"9fe0800c",
   936 => x"0294050d",
   937 => x"0402cc05",
   938 => x"0d7e605e",
   939 => x"5b8056ff",
   940 => x"0b9fe5d8",
   941 => x"0c9fe1c0",
   942 => x"089fe5e4",
   943 => x"0856579f",
   944 => x"e5ec0876",
   945 => x"2e8e389f",
   946 => x"e5f40884",
   947 => x"2b598480",
   948 => x"809ddb04",
   949 => x"9fe5f008",
   950 => x"842b5980",
   951 => x"5a797927",
   952 => x"81e83879",
   953 => x"8f06a017",
   954 => x"575473a2",
   955 => x"38745284",
   956 => x"8080a6d0",
   957 => x"51848080",
   958 => x"82832d9f",
   959 => x"e1c45274",
   960 => x"51811555",
   961 => x"84808090",
   962 => x"d72d9fe1",
   963 => x"c4568076",
   964 => x"84808080",
   965 => x"f52d5558",
   966 => x"73782e83",
   967 => x"38815873",
   968 => x"81e52e81",
   969 => x"9c388170",
   970 => x"7906555c",
   971 => x"73802e81",
   972 => x"90388b16",
   973 => x"84808080",
   974 => x"f52d9806",
   975 => x"58778181",
   976 => x"388b537c",
   977 => x"52755184",
   978 => x"808093df",
   979 => x"2d9fe080",
   980 => x"0880ee38",
   981 => x"9c160851",
   982 => x"84808084",
   983 => x"eb2d9fe0",
   984 => x"8008841c",
   985 => x"0c9a1684",
   986 => x"808080e0",
   987 => x"2d518480",
   988 => x"80859c2d",
   989 => x"9fe08008",
   990 => x"9fe08008",
   991 => x"55559fe5",
   992 => x"ec08802e",
   993 => x"9f389416",
   994 => x"84808080",
   995 => x"e02d5184",
   996 => x"8080859c",
   997 => x"2d9fe080",
   998 => x"08902b83",
   999 => x"fff00a06",
  1000 => x"70165154",
  1001 => x"73881c0c",
  1002 => x"777b0c7c",
  1003 => x"52848080",
  1004 => x"a6f05184",
  1005 => x"80808283",
  1006 => x"2d7b5484",
  1007 => x"8080a097",
  1008 => x"04811a5a",
  1009 => x"8480809d",
  1010 => x"dd049fe5",
  1011 => x"ec08802e",
  1012 => x"80c33876",
  1013 => x"51848080",
  1014 => x"9c8f2d9f",
  1015 => x"e080089f",
  1016 => x"e0800853",
  1017 => x"848080a7",
  1018 => x"84525784",
  1019 => x"80808283",
  1020 => x"2d7680ff",
  1021 => x"fffff806",
  1022 => x"547380ff",
  1023 => x"fffff82e",
  1024 => x"9438fe17",
  1025 => x"9fe5f408",
  1026 => x"299fe5fc",
  1027 => x"08055584",
  1028 => x"80809ddb",
  1029 => x"04805473",
  1030 => x"9fe0800c",
  1031 => x"02b4050d",
  1032 => x"0402e405",
  1033 => x"0d787a71",
  1034 => x"549fe5c8",
  1035 => x"53555584",
  1036 => x"80809da5",
  1037 => x"2d9fe080",
  1038 => x"0881ff06",
  1039 => x"5372802e",
  1040 => x"80fe3884",
  1041 => x"8080a79c",
  1042 => x"51848080",
  1043 => x"92b12d9f",
  1044 => x"e5cc0883",
  1045 => x"ff05892a",
  1046 => x"57807056",
  1047 => x"56757725",
  1048 => x"80fd389f",
  1049 => x"e5d008fe",
  1050 => x"059fe5f4",
  1051 => x"08299fe5",
  1052 => x"fc081176",
  1053 => x"9fe5e808",
  1054 => x"06057554",
  1055 => x"52538480",
  1056 => x"8090d72d",
  1057 => x"9fe08008",
  1058 => x"802e80c8",
  1059 => x"38811570",
  1060 => x"9fe5e808",
  1061 => x"06545572",
  1062 => x"94389fe5",
  1063 => x"d0085184",
  1064 => x"80809c8f",
  1065 => x"2d9fe080",
  1066 => x"089fe5d0",
  1067 => x"0c848014",
  1068 => x"81175754",
  1069 => x"767624ff",
  1070 => x"aa388480",
  1071 => x"80a1df04",
  1072 => x"74528480",
  1073 => x"80a7b851",
  1074 => x"84808082",
  1075 => x"832d8480",
  1076 => x"80a1e104",
  1077 => x"9fe08008",
  1078 => x"53848080",
  1079 => x"a1e10481",
  1080 => x"53729fe0",
  1081 => x"800c029c",
  1082 => x"050d0400",
  1083 => x"00ffffff",
  1084 => x"ff00ffff",
  1085 => x"ffff00ff",
  1086 => x"ffffff00",
  1087 => x"476f7420",
  1088 => x"72657375",
  1089 => x"6c742025",
  1090 => x"64200a00",
  1091 => x"434d4435",
  1092 => x"35202564",
  1093 => x"0a000000",
  1094 => x"434d4434",
  1095 => x"31202564",
  1096 => x"0a000000",
  1097 => x"436d645f",
  1098 => x"696e6974",
  1099 => x"0a000000",
  1100 => x"696e6974",
  1101 => x"2025640a",
  1102 => x"20200000",
  1103 => x"636d645f",
  1104 => x"434d4438",
  1105 => x"20726573",
  1106 => x"706f6e73",
  1107 => x"653a2025",
  1108 => x"640a0000",
  1109 => x"434d4438",
  1110 => x"5f342072",
  1111 => x"6573706f",
  1112 => x"6e73653a",
  1113 => x"2025640a",
  1114 => x"00000000",
  1115 => x"53444843",
  1116 => x"20496e69",
  1117 => x"7469616c",
  1118 => x"697a6174",
  1119 => x"696f6e20",
  1120 => x"6572726f",
  1121 => x"72210a00",
  1122 => x"434d4435",
  1123 => x"38202564",
  1124 => x"0a202000",
  1125 => x"434d4435",
  1126 => x"385f3220",
  1127 => x"25640a20",
  1128 => x"20000000",
  1129 => x"73645f72",
  1130 => x"6561645f",
  1131 => x"73656374",
  1132 => x"6f722025",
  1133 => x"642c2025",
  1134 => x"640a0000",
  1135 => x"52656164",
  1136 => x"20636f6d",
  1137 => x"6d616e64",
  1138 => x"20666169",
  1139 => x"6c656420",
  1140 => x"61742025",
  1141 => x"64202825",
  1142 => x"64290a00",
  1143 => x"496e6974",
  1144 => x"69616c69",
  1145 => x"7a696e67",
  1146 => x"20534420",
  1147 => x"63617264",
  1148 => x"0a000000",
  1149 => x"48756e74",
  1150 => x"696e6720",
  1151 => x"666f7220",
  1152 => x"70617274",
  1153 => x"6974696f",
  1154 => x"6e0a0000",
  1155 => x"4f53445a",
  1156 => x"50553031",
  1157 => x"53595300",
  1158 => x"43616e27",
  1159 => x"74206c6f",
  1160 => x"61642066",
  1161 => x"69726d77",
  1162 => x"6172650a",
  1163 => x"00000000",
  1164 => x"4661696c",
  1165 => x"65642074",
  1166 => x"6f20696e",
  1167 => x"69746961",
  1168 => x"6c697a65",
  1169 => x"20534420",
  1170 => x"63617264",
  1171 => x"0a000000",
  1172 => x"52656164",
  1173 => x"696e6720",
  1174 => x"4d42520a",
  1175 => x"00000000",
  1176 => x"52656164",
  1177 => x"206f6620",
  1178 => x"4d425220",
  1179 => x"6661696c",
  1180 => x"65640a00",
  1181 => x"4d425220",
  1182 => x"73756363",
  1183 => x"65737366",
  1184 => x"756c6c79",
  1185 => x"20726561",
  1186 => x"640a0000",
  1187 => x"46415431",
  1188 => x"36202020",
  1189 => x"00000000",
  1190 => x"46415433",
  1191 => x"32202020",
  1192 => x"00000000",
  1193 => x"50617274",
  1194 => x"6974696f",
  1195 => x"6e636f75",
  1196 => x"6e742025",
  1197 => x"640a0000",
  1198 => x"4e6f2070",
  1199 => x"61727469",
  1200 => x"74696f6e",
  1201 => x"20736967",
  1202 => x"6e617475",
  1203 => x"72652066",
  1204 => x"6f756e64",
  1205 => x"0a000000",
  1206 => x"52656164",
  1207 => x"696e6720",
  1208 => x"626f6f74",
  1209 => x"20736563",
  1210 => x"746f7220",
  1211 => x"25640a00",
  1212 => x"52656164",
  1213 => x"20626f6f",
  1214 => x"74207365",
  1215 => x"63746f72",
  1216 => x"2066726f",
  1217 => x"6d206669",
  1218 => x"72737420",
  1219 => x"70617274",
  1220 => x"6974696f",
  1221 => x"6e0a0000",
  1222 => x"48756e74",
  1223 => x"696e6720",
  1224 => x"666f7220",
  1225 => x"66696c65",
  1226 => x"73797374",
  1227 => x"656d0a00",
  1228 => x"556e7375",
  1229 => x"70706f72",
  1230 => x"74656420",
  1231 => x"70617274",
  1232 => x"6974696f",
  1233 => x"6e207479",
  1234 => x"7065210d",
  1235 => x"00000000",
  1236 => x"52656164",
  1237 => x"696e6720",
  1238 => x"64697265",
  1239 => x"63746f72",
  1240 => x"79207365",
  1241 => x"63746f72",
  1242 => x"2025640a",
  1243 => x"00000000",
  1244 => x"66696c65",
  1245 => x"20222573",
  1246 => x"2220666f",
  1247 => x"756e640d",
  1248 => x"00000000",
  1249 => x"47657446",
  1250 => x"41544c69",
  1251 => x"6e6b2072",
  1252 => x"65747572",
  1253 => x"6e656420",
  1254 => x"25640a00",
  1255 => x"4f70656e",
  1256 => x"65642066",
  1257 => x"696c652c",
  1258 => x"206c6f61",
  1259 => x"64696e67",
  1260 => x"2e2e2e0a",
  1261 => x"00000000",
  1262 => x"43616e27",
  1263 => x"74206f70",
  1264 => x"656e2025",
  1265 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

