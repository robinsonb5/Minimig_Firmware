library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity amigaboot_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM downto 0);
	q : out std_logic_vector(15 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(15 downto 0) := X"0000";
	we_n : in std_logic := '1';
	uds_n : in std_logic := '1';
	lds_n : in std_logic := '1'
);
end amigaboot_ROM;

architecture arch of amigaboot_ROM is

type ram_type is array(natural range 0 to (2**(maxAddrBitBRAM+1)-1)) of std_logic_vector(7 downto 0);

shared variable ram : ram_type :=
(
     0 => x"00",
     1 => x"01",
     2 => x"00",
     3 => x"00",
     4 => x"00",
     5 => x"00",
     6 => x"00",
     7 => x"08",
     8 => x"4d",
     9 => x"f9",
    10 => x"00",
    11 => x"df",
    12 => x"f0",
    13 => x"00",
    14 => x"3d",
    15 => x"7c",
    16 => x"90",
    17 => x"00",
    18 => x"01",
    19 => x"00",
    20 => x"3d",
    21 => x"7c",
    22 => x"00",
    23 => x"00",
    24 => x"01",
    25 => x"02",
    26 => x"3d",
    27 => x"7c",
    28 => x"00",
    29 => x"00",
    30 => x"01",
    31 => x"04",
    32 => x"3d",
    33 => x"7c",
    34 => x"00",
    35 => x"00",
    36 => x"01",
    37 => x"08",
    38 => x"3d",
    39 => x"7c",
    40 => x"00",
    41 => x"00",
    42 => x"01",
    43 => x"0a",
    44 => x"61",
    45 => x"00",
    46 => x"02",
    47 => x"de",
    48 => x"3d",
    49 => x"7c",
    50 => x"00",
    51 => x"3c",
    52 => x"00",
    53 => x"92",
    54 => x"3d",
    55 => x"7c",
    56 => x"00",
    57 => x"d4",
    58 => x"00",
    59 => x"94",
    60 => x"3d",
    61 => x"7c",
    62 => x"2c",
    63 => x"81",
    64 => x"00",
    65 => x"8e",
    66 => x"3d",
    67 => x"7c",
    68 => x"f4",
    69 => x"c1",
    70 => x"00",
    71 => x"90",
    72 => x"3d",
    73 => x"7c",
    74 => x"03",
    75 => x"7f",
    76 => x"01",
    77 => x"80",
    78 => x"3d",
    79 => x"7c",
    80 => x"0f",
    81 => x"ff",
    82 => x"01",
    83 => x"82",
    84 => x"41",
    85 => x"fa",
    86 => x"02",
    87 => x"d2",
    88 => x"43",
    89 => x"f9",
    90 => x"00",
    91 => x"00",
    92 => x"c1",
    93 => x"00",
    94 => x"70",
    95 => x"02",
    96 => x"22",
    97 => x"d8",
    98 => x"4e",
    99 => x"71",
   100 => x"51",
   101 => x"c8",
   102 => x"ff",
   103 => x"fa",
   104 => x"2d",
   105 => x"7c",
   106 => x"00",
   107 => x"00",
   108 => x"c1",
   109 => x"00",
   110 => x"00",
   111 => x"80",
   112 => x"3d",
   113 => x"40",
   114 => x"00",
   115 => x"88",
   116 => x"3d",
   117 => x"7c",
   118 => x"83",
   119 => x"90",
   120 => x"00",
   121 => x"96",
   122 => x"3d",
   123 => x"7c",
   124 => x"7f",
   125 => x"ff",
   126 => x"00",
   127 => x"9e",
   128 => x"41",
   129 => x"fa",
   130 => x"06",
   131 => x"4b",
   132 => x"61",
   133 => x"00",
   134 => x"02",
   135 => x"5e",
   136 => x"41",
   137 => x"fa",
   138 => x"06",
   139 => x"e3",
   140 => x"61",
   141 => x"00",
   142 => x"02",
   143 => x"56",
   144 => x"41",
   145 => x"fa",
   146 => x"06",
   147 => x"f5",
   148 => x"61",
   149 => x"00",
   150 => x"02",
   151 => x"4e",
   152 => x"41",
   153 => x"fa",
   154 => x"05",
   155 => x"9a",
   156 => x"61",
   157 => x"00",
   158 => x"02",
   159 => x"46",
   160 => x"30",
   161 => x"2e",
   162 => x"00",
   163 => x"04",
   164 => x"e0",
   165 => x"48",
   166 => x"02",
   167 => x"00",
   168 => x"00",
   169 => x"7f",
   170 => x"61",
   171 => x"00",
   172 => x"01",
   173 => x"d0",
   174 => x"41",
   175 => x"fa",
   176 => x"05",
   177 => x"92",
   178 => x"08",
   179 => x"01",
   180 => x"00",
   181 => x"04",
   182 => x"67",
   183 => x"04",
   184 => x"41",
   185 => x"fa",
   186 => x"05",
   187 => x"8f",
   188 => x"61",
   189 => x"00",
   190 => x"02",
   191 => x"26",
   192 => x"41",
   193 => x"fa",
   194 => x"05",
   195 => x"8f",
   196 => x"61",
   197 => x"00",
   198 => x"02",
   199 => x"1e",
   200 => x"30",
   201 => x"2e",
   202 => x"00",
   203 => x"7c",
   204 => x"61",
   205 => x"00",
   206 => x"01",
   207 => x"ae",
   208 => x"70",
   209 => x"0a",
   210 => x"61",
   211 => x"00",
   212 => x"01",
   213 => x"c0",
   214 => x"70",
   215 => x"0a",
   216 => x"61",
   217 => x"00",
   218 => x"01",
   219 => x"ba",
   220 => x"13",
   221 => x"fc",
   222 => x"00",
   223 => x"03",
   224 => x"00",
   225 => x"bf",
   226 => x"e2",
   227 => x"01",
   228 => x"13",
   229 => x"fc",
   230 => x"00",
   231 => x"00",
   232 => x"00",
   233 => x"bf",
   234 => x"e0",
   235 => x"01",
   236 => x"13",
   237 => x"fc",
   238 => x"00",
   239 => x"ff",
   240 => x"00",
   241 => x"bf",
   242 => x"d3",
   243 => x"00",
   244 => x"13",
   245 => x"fc",
   246 => x"00",
   247 => x"f7",
   248 => x"00",
   249 => x"bf",
   250 => x"d1",
   251 => x"00",
   252 => x"13",
   253 => x"fc",
   254 => x"00",
   255 => x"f6",
   256 => x"00",
   257 => x"bf",
   258 => x"d1",
   259 => x"00",
   260 => x"13",
   261 => x"fc",
   262 => x"00",
   263 => x"f7",
   264 => x"00",
   265 => x"bf",
   266 => x"d1",
   267 => x"00",
   268 => x"08",
   269 => x"39",
   270 => x"00",
   271 => x"02",
   272 => x"00",
   273 => x"bf",
   274 => x"e0",
   275 => x"01",
   276 => x"67",
   277 => x"e6",
   278 => x"30",
   279 => x"3c",
   280 => x"00",
   281 => x"0c",
   282 => x"61",
   283 => x"00",
   284 => x"01",
   285 => x"28",
   286 => x"30",
   287 => x"7c",
   288 => x"40",
   289 => x"00",
   290 => x"0c",
   291 => x"58",
   292 => x"aa",
   293 => x"ca",
   294 => x"66",
   295 => x"00",
   296 => x"01",
   297 => x"08",
   298 => x"30",
   299 => x"18",
   300 => x"b0",
   301 => x"7c",
   302 => x"00",
   303 => x"01",
   304 => x"66",
   305 => x"26",
   306 => x"20",
   307 => x"18",
   308 => x"61",
   309 => x"00",
   310 => x"01",
   311 => x"0e",
   312 => x"41",
   313 => x"f8",
   314 => x"40",
   315 => x"00",
   316 => x"0c",
   317 => x"10",
   318 => x"00",
   319 => x"fe",
   320 => x"66",
   321 => x"08",
   322 => x"3d",
   323 => x"7c",
   324 => x"0f",
   325 => x"00",
   326 => x"01",
   327 => x"80",
   328 => x"52",
   329 => x"48",
   330 => x"61",
   331 => x"00",
   332 => x"01",
   333 => x"98",
   334 => x"70",
   335 => x"0a",
   336 => x"61",
   337 => x"00",
   338 => x"01",
   339 => x"42",
   340 => x"60",
   341 => x"00",
   342 => x"00",
   343 => x"ea",
   344 => x"b0",
   345 => x"7c",
   346 => x"00",
   347 => x"02",
   348 => x"66",
   349 => x"00",
   350 => x"00",
   351 => x"92",
   352 => x"28",
   353 => x"58",
   354 => x"2a",
   355 => x"4c",
   356 => x"28",
   357 => x"18",
   358 => x"2a",
   359 => x"04",
   360 => x"41",
   361 => x"fa",
   362 => x"04",
   363 => x"f5",
   364 => x"61",
   365 => x"00",
   366 => x"01",
   367 => x"76",
   368 => x"20",
   369 => x"0c",
   370 => x"61",
   371 => x"00",
   372 => x"00",
   373 => x"f8",
   374 => x"41",
   375 => x"fa",
   376 => x"04",
   377 => x"f6",
   378 => x"61",
   379 => x"00",
   380 => x"01",
   381 => x"68",
   382 => x"20",
   383 => x"04",
   384 => x"61",
   385 => x"00",
   386 => x"00",
   387 => x"ea",
   388 => x"70",
   389 => x"0a",
   390 => x"61",
   391 => x"00",
   392 => x"01",
   393 => x"0c",
   394 => x"41",
   395 => x"fa",
   396 => x"04",
   397 => x"ec",
   398 => x"61",
   399 => x"00",
   400 => x"01",
   401 => x"54",
   402 => x"94",
   403 => x"7c",
   404 => x"00",
   405 => x"21",
   406 => x"47",
   407 => x"eb",
   408 => x"ff",
   409 => x"df",
   410 => x"2c",
   411 => x"05",
   412 => x"ea",
   413 => x"8e",
   414 => x"bc",
   415 => x"84",
   416 => x"6d",
   417 => x"02",
   418 => x"2c",
   419 => x"04",
   420 => x"30",
   421 => x"06",
   422 => x"61",
   423 => x"00",
   424 => x"00",
   425 => x"9c",
   426 => x"30",
   427 => x"06",
   428 => x"e4",
   429 => x"48",
   430 => x"53",
   431 => x"40",
   432 => x"28",
   433 => x"d8",
   434 => x"4e",
   435 => x"71",
   436 => x"51",
   437 => x"c8",
   438 => x"ff",
   439 => x"fa",
   440 => x"70",
   441 => x"7f",
   442 => x"61",
   443 => x"00",
   444 => x"00",
   445 => x"d8",
   446 => x"08",
   447 => x"79",
   448 => x"00",
   449 => x"01",
   450 => x"00",
   451 => x"bf",
   452 => x"e0",
   453 => x"01",
   454 => x"98",
   455 => x"86",
   456 => x"6e",
   457 => x"d0",
   458 => x"bb",
   459 => x"fc",
   460 => x"00",
   461 => x"f8",
   462 => x"00",
   463 => x"00",
   464 => x"66",
   465 => x"16",
   466 => x"ba",
   467 => x"bc",
   468 => x"00",
   469 => x"04",
   470 => x"00",
   471 => x"00",
   472 => x"66",
   473 => x"0e",
   474 => x"28",
   475 => x"4d",
   476 => x"d9",
   477 => x"c5",
   478 => x"7a",
   479 => x"ff",
   480 => x"28",
   481 => x"dd",
   482 => x"4e",
   483 => x"71",
   484 => x"51",
   485 => x"cd",
   486 => x"ff",
   487 => x"fa",
   488 => x"70",
   489 => x"0a",
   490 => x"61",
   491 => x"00",
   492 => x"00",
   493 => x"a8",
   494 => x"60",
   495 => x"50",
   496 => x"b0",
   497 => x"7c",
   498 => x"00",
   499 => x"03",
   500 => x"66",
   501 => x"10",
   502 => x"08",
   503 => x"f9",
   504 => x"00",
   505 => x"01",
   506 => x"00",
   507 => x"bf",
   508 => x"e0",
   509 => x"01",
   510 => x"4a",
   511 => x"39",
   512 => x"00",
   513 => x"bf",
   514 => x"c0",
   515 => x"00",
   516 => x"60",
   517 => x"fe",
   518 => x"b0",
   519 => x"7c",
   520 => x"00",
   521 => x"04",
   522 => x"66",
   523 => x"0e",
   524 => x"28",
   525 => x"58",
   526 => x"28",
   527 => x"18",
   528 => x"70",
   529 => x"00",
   530 => x"28",
   531 => x"c0",
   532 => x"59",
   533 => x"84",
   534 => x"6e",
   535 => x"fa",
   536 => x"60",
   537 => x"26",
   538 => x"3e",
   539 => x"00",
   540 => x"3d",
   541 => x"7c",
   542 => x"0f",
   543 => x"00",
   544 => x"01",
   545 => x"80",
   546 => x"41",
   547 => x"fa",
   548 => x"04",
   549 => x"95",
   550 => x"61",
   551 => x"00",
   552 => x"00",
   553 => x"bc",
   554 => x"30",
   555 => x"07",
   556 => x"61",
   557 => x"46",
   558 => x"60",
   559 => x"fe",
   560 => x"3d",
   561 => x"7c",
   562 => x"0f",
   563 => x"00",
   564 => x"01",
   565 => x"80",
   566 => x"41",
   567 => x"fa",
   568 => x"04",
   569 => x"63",
   570 => x"61",
   571 => x"00",
   572 => x"00",
   573 => x"a8",
   574 => x"60",
   575 => x"ee",
   576 => x"60",
   577 => x"00",
   578 => x"fe",
   579 => x"d4",
   580 => x"3d",
   581 => x"7c",
   582 => x"00",
   583 => x"02",
   584 => x"00",
   585 => x"9c",
   586 => x"30",
   587 => x"7c",
   588 => x"40",
   589 => x"00",
   590 => x"2d",
   591 => x"48",
   592 => x"00",
   593 => x"20",
   594 => x"e2",
   595 => x"48",
   596 => x"00",
   597 => x"40",
   598 => x"80",
   599 => x"00",
   600 => x"3d",
   601 => x"40",
   602 => x"00",
   603 => x"24",
   604 => x"3d",
   605 => x"40",
   606 => x"00",
   607 => x"24",
   608 => x"30",
   609 => x"2e",
   610 => x"00",
   611 => x"1e",
   612 => x"08",
   613 => x"00",
   614 => x"00",
   615 => x"01",
   616 => x"67",
   617 => x"f6",
   618 => x"4e",
   619 => x"75",
   620 => x"48",
   621 => x"40",
   622 => x"61",
   623 => x"04",
   624 => x"48",
   625 => x"41",
   626 => x"20",
   627 => x"01",
   628 => x"e0",
   629 => x"58",
   630 => x"61",
   631 => x"04",
   632 => x"20",
   633 => x"01",
   634 => x"e0",
   635 => x"58",
   636 => x"22",
   637 => x"00",
   638 => x"e8",
   639 => x"08",
   640 => x"61",
   641 => x"06",
   642 => x"20",
   643 => x"01",
   644 => x"02",
   645 => x"00",
   646 => x"00",
   647 => x"0f",
   648 => x"d0",
   649 => x"3c",
   650 => x"00",
   651 => x"30",
   652 => x"b0",
   653 => x"3c",
   654 => x"00",
   655 => x"39",
   656 => x"6f",
   657 => x"02",
   658 => x"5e",
   659 => x"00",
   660 => x"22",
   661 => x"4b",
   662 => x"52",
   663 => x"8b",
   664 => x"b0",
   665 => x"3c",
   666 => x"00",
   667 => x"0a",
   668 => x"66",
   669 => x"0c",
   670 => x"96",
   671 => x"c2",
   672 => x"34",
   673 => x"3c",
   674 => x"00",
   675 => x"00",
   676 => x"47",
   677 => x"eb",
   678 => x"02",
   679 => x"7f",
   680 => x"60",
   681 => x"28",
   682 => x"48",
   683 => x"80",
   684 => x"90",
   685 => x"7c",
   686 => x"00",
   687 => x"20",
   688 => x"e7",
   689 => x"40",
   690 => x"41",
   691 => x"fa",
   692 => x"00",
   693 => x"80",
   694 => x"d0",
   695 => x"c0",
   696 => x"70",
   697 => x"07",
   698 => x"12",
   699 => x"98",
   700 => x"43",
   701 => x"e9",
   702 => x"00",
   703 => x"50",
   704 => x"51",
   705 => x"c8",
   706 => x"ff",
   707 => x"f8",
   708 => x"52",
   709 => x"42",
   710 => x"b4",
   711 => x"7c",
   712 => x"00",
   713 => x"50",
   714 => x"66",
   715 => x"16",
   716 => x"74",
   717 => x"00",
   718 => x"47",
   719 => x"eb",
   720 => x"02",
   721 => x"30",
   722 => x"52",
   723 => x"43",
   724 => x"b6",
   725 => x"7c",
   726 => x"00",
   727 => x"19",
   728 => x"66",
   729 => x"08",
   730 => x"53",
   731 => x"43",
   732 => x"47",
   733 => x"eb",
   734 => x"fd",
   735 => x"80",
   736 => x"61",
   737 => x"12",
   738 => x"4e",
   739 => x"75",
   740 => x"24",
   741 => x"48",
   742 => x"22",
   743 => x"4b",
   744 => x"70",
   745 => x"00",
   746 => x"10",
   747 => x"1a",
   748 => x"67",
   749 => x"04",
   750 => x"61",
   751 => x"a4",
   752 => x"60",
   753 => x"f4",
   754 => x"4e",
   755 => x"75",
   756 => x"41",
   757 => x"f9",
   758 => x"00",
   759 => x"00",
   760 => x"80",
   761 => x"00",
   762 => x"43",
   763 => x"e8",
   764 => x"02",
   765 => x"80",
   766 => x"30",
   767 => x"3c",
   768 => x"0f",
   769 => x"9f",
   770 => x"20",
   771 => x"d9",
   772 => x"4e",
   773 => x"71",
   774 => x"51",
   775 => x"c8",
   776 => x"ff",
   777 => x"fa",
   778 => x"4e",
   779 => x"75",
   780 => x"74",
   781 => x"00",
   782 => x"76",
   783 => x"00",
   784 => x"47",
   785 => x"f9",
   786 => x"00",
   787 => x"00",
   788 => x"80",
   789 => x"00",
   790 => x"20",
   791 => x"4b",
   792 => x"70",
   793 => x"00",
   794 => x"32",
   795 => x"3c",
   796 => x"10",
   797 => x"3f",
   798 => x"20",
   799 => x"c0",
   800 => x"4e",
   801 => x"71",
   802 => x"51",
   803 => x"c9",
   804 => x"ff",
   805 => x"fa",
   806 => x"4e",
   807 => x"75",
   808 => x"00",
   809 => x"e0",
   810 => x"00",
   811 => x"00",
   812 => x"00",
   813 => x"e2",
   814 => x"80",
   815 => x"00",
   816 => x"ff",
   817 => x"ff",
   818 => x"ff",
   819 => x"fe",
   820 => x"00",
   821 => x"00",
   822 => x"00",
   823 => x"00",
   824 => x"00",
   825 => x"00",
   826 => x"00",
   827 => x"00",
   828 => x"18",
   829 => x"18",
   830 => x"18",
   831 => x"18",
   832 => x"18",
   833 => x"00",
   834 => x"18",
   835 => x"00",
   836 => x"6c",
   837 => x"6c",
   838 => x"00",
   839 => x"00",
   840 => x"00",
   841 => x"00",
   842 => x"00",
   843 => x"00",
   844 => x"6c",
   845 => x"6c",
   846 => x"fe",
   847 => x"6c",
   848 => x"fe",
   849 => x"6c",
   850 => x"6c",
   851 => x"00",
   852 => x"18",
   853 => x"3e",
   854 => x"60",
   855 => x"3c",
   856 => x"06",
   857 => x"7c",
   858 => x"18",
   859 => x"00",
   860 => x"00",
   861 => x"66",
   862 => x"ac",
   863 => x"d8",
   864 => x"36",
   865 => x"6a",
   866 => x"cc",
   867 => x"00",
   868 => x"38",
   869 => x"6c",
   870 => x"68",
   871 => x"76",
   872 => x"dc",
   873 => x"ce",
   874 => x"7b",
   875 => x"00",
   876 => x"18",
   877 => x"18",
   878 => x"30",
   879 => x"00",
   880 => x"00",
   881 => x"00",
   882 => x"00",
   883 => x"00",
   884 => x"0c",
   885 => x"18",
   886 => x"30",
   887 => x"30",
   888 => x"30",
   889 => x"18",
   890 => x"0c",
   891 => x"00",
   892 => x"30",
   893 => x"18",
   894 => x"0c",
   895 => x"0c",
   896 => x"0c",
   897 => x"18",
   898 => x"30",
   899 => x"00",
   900 => x"00",
   901 => x"66",
   902 => x"3c",
   903 => x"ff",
   904 => x"3c",
   905 => x"66",
   906 => x"00",
   907 => x"00",
   908 => x"00",
   909 => x"18",
   910 => x"18",
   911 => x"7e",
   912 => x"18",
   913 => x"18",
   914 => x"00",
   915 => x"00",
   916 => x"00",
   917 => x"00",
   918 => x"00",
   919 => x"00",
   920 => x"00",
   921 => x"18",
   922 => x"18",
   923 => x"30",
   924 => x"00",
   925 => x"00",
   926 => x"00",
   927 => x"7e",
   928 => x"00",
   929 => x"00",
   930 => x"00",
   931 => x"00",
   932 => x"00",
   933 => x"00",
   934 => x"00",
   935 => x"00",
   936 => x"00",
   937 => x"18",
   938 => x"18",
   939 => x"00",
   940 => x"03",
   941 => x"06",
   942 => x"0c",
   943 => x"18",
   944 => x"30",
   945 => x"60",
   946 => x"c0",
   947 => x"00",
   948 => x"3c",
   949 => x"66",
   950 => x"6e",
   951 => x"7e",
   952 => x"76",
   953 => x"66",
   954 => x"3c",
   955 => x"00",
   956 => x"18",
   957 => x"38",
   958 => x"78",
   959 => x"18",
   960 => x"18",
   961 => x"18",
   962 => x"18",
   963 => x"00",
   964 => x"3c",
   965 => x"66",
   966 => x"06",
   967 => x"0c",
   968 => x"18",
   969 => x"30",
   970 => x"7e",
   971 => x"00",
   972 => x"3c",
   973 => x"66",
   974 => x"06",
   975 => x"1c",
   976 => x"06",
   977 => x"66",
   978 => x"3c",
   979 => x"00",
   980 => x"1c",
   981 => x"3c",
   982 => x"6c",
   983 => x"cc",
   984 => x"fe",
   985 => x"0c",
   986 => x"0c",
   987 => x"00",
   988 => x"7e",
   989 => x"60",
   990 => x"7c",
   991 => x"06",
   992 => x"06",
   993 => x"66",
   994 => x"3c",
   995 => x"00",
   996 => x"1c",
   997 => x"30",
   998 => x"60",
   999 => x"7c",
  1000 => x"66",
  1001 => x"66",
  1002 => x"3c",
  1003 => x"00",
  1004 => x"7e",
  1005 => x"06",
  1006 => x"06",
  1007 => x"0c",
  1008 => x"18",
  1009 => x"18",
  1010 => x"18",
  1011 => x"00",
  1012 => x"3c",
  1013 => x"66",
  1014 => x"66",
  1015 => x"3c",
  1016 => x"66",
  1017 => x"66",
  1018 => x"3c",
  1019 => x"00",
  1020 => x"3c",
  1021 => x"66",
  1022 => x"66",
  1023 => x"3e",
  1024 => x"06",
  1025 => x"0c",
  1026 => x"38",
  1027 => x"00",
  1028 => x"00",
  1029 => x"18",
  1030 => x"18",
  1031 => x"00",
  1032 => x"00",
  1033 => x"18",
  1034 => x"18",
  1035 => x"00",
  1036 => x"00",
  1037 => x"18",
  1038 => x"18",
  1039 => x"00",
  1040 => x"00",
  1041 => x"18",
  1042 => x"18",
  1043 => x"30",
  1044 => x"00",
  1045 => x"06",
  1046 => x"18",
  1047 => x"60",
  1048 => x"18",
  1049 => x"06",
  1050 => x"00",
  1051 => x"00",
  1052 => x"00",
  1053 => x"00",
  1054 => x"7e",
  1055 => x"00",
  1056 => x"7e",
  1057 => x"00",
  1058 => x"00",
  1059 => x"00",
  1060 => x"00",
  1061 => x"60",
  1062 => x"18",
  1063 => x"06",
  1064 => x"18",
  1065 => x"60",
  1066 => x"00",
  1067 => x"00",
  1068 => x"3c",
  1069 => x"66",
  1070 => x"06",
  1071 => x"0c",
  1072 => x"18",
  1073 => x"00",
  1074 => x"18",
  1075 => x"00",
  1076 => x"7c",
  1077 => x"c6",
  1078 => x"de",
  1079 => x"d6",
  1080 => x"de",
  1081 => x"c0",
  1082 => x"78",
  1083 => x"00",
  1084 => x"3c",
  1085 => x"66",
  1086 => x"66",
  1087 => x"7e",
  1088 => x"66",
  1089 => x"66",
  1090 => x"66",
  1091 => x"00",
  1092 => x"7c",
  1093 => x"66",
  1094 => x"66",
  1095 => x"7c",
  1096 => x"66",
  1097 => x"66",
  1098 => x"7c",
  1099 => x"00",
  1100 => x"1e",
  1101 => x"30",
  1102 => x"60",
  1103 => x"60",
  1104 => x"60",
  1105 => x"30",
  1106 => x"1e",
  1107 => x"00",
  1108 => x"78",
  1109 => x"6c",
  1110 => x"66",
  1111 => x"66",
  1112 => x"66",
  1113 => x"6c",
  1114 => x"78",
  1115 => x"00",
  1116 => x"7e",
  1117 => x"60",
  1118 => x"60",
  1119 => x"78",
  1120 => x"60",
  1121 => x"60",
  1122 => x"7e",
  1123 => x"00",
  1124 => x"7e",
  1125 => x"60",
  1126 => x"60",
  1127 => x"78",
  1128 => x"60",
  1129 => x"60",
  1130 => x"60",
  1131 => x"00",
  1132 => x"3c",
  1133 => x"66",
  1134 => x"60",
  1135 => x"6e",
  1136 => x"66",
  1137 => x"66",
  1138 => x"3e",
  1139 => x"00",
  1140 => x"66",
  1141 => x"66",
  1142 => x"66",
  1143 => x"7e",
  1144 => x"66",
  1145 => x"66",
  1146 => x"66",
  1147 => x"00",
  1148 => x"3c",
  1149 => x"18",
  1150 => x"18",
  1151 => x"18",
  1152 => x"18",
  1153 => x"18",
  1154 => x"3c",
  1155 => x"00",
  1156 => x"06",
  1157 => x"06",
  1158 => x"06",
  1159 => x"06",
  1160 => x"06",
  1161 => x"66",
  1162 => x"3c",
  1163 => x"00",
  1164 => x"c6",
  1165 => x"cc",
  1166 => x"d8",
  1167 => x"f0",
  1168 => x"d8",
  1169 => x"cc",
  1170 => x"c6",
  1171 => x"00",
  1172 => x"60",
  1173 => x"60",
  1174 => x"60",
  1175 => x"60",
  1176 => x"60",
  1177 => x"60",
  1178 => x"7e",
  1179 => x"00",
  1180 => x"c6",
  1181 => x"ee",
  1182 => x"fe",
  1183 => x"d6",
  1184 => x"c6",
  1185 => x"c6",
  1186 => x"c6",
  1187 => x"00",
  1188 => x"c6",
  1189 => x"e6",
  1190 => x"f6",
  1191 => x"de",
  1192 => x"ce",
  1193 => x"c6",
  1194 => x"c6",
  1195 => x"00",
  1196 => x"3c",
  1197 => x"66",
  1198 => x"66",
  1199 => x"66",
  1200 => x"66",
  1201 => x"66",
  1202 => x"3c",
  1203 => x"00",
  1204 => x"7c",
  1205 => x"66",
  1206 => x"66",
  1207 => x"7c",
  1208 => x"60",
  1209 => x"60",
  1210 => x"60",
  1211 => x"00",
  1212 => x"78",
  1213 => x"cc",
  1214 => x"cc",
  1215 => x"cc",
  1216 => x"cc",
  1217 => x"dc",
  1218 => x"7e",
  1219 => x"00",
  1220 => x"7c",
  1221 => x"66",
  1222 => x"66",
  1223 => x"7c",
  1224 => x"6c",
  1225 => x"66",
  1226 => x"66",
  1227 => x"00",
  1228 => x"3c",
  1229 => x"66",
  1230 => x"70",
  1231 => x"3c",
  1232 => x"0e",
  1233 => x"66",
  1234 => x"3c",
  1235 => x"00",
  1236 => x"7e",
  1237 => x"18",
  1238 => x"18",
  1239 => x"18",
  1240 => x"18",
  1241 => x"18",
  1242 => x"18",
  1243 => x"00",
  1244 => x"66",
  1245 => x"66",
  1246 => x"66",
  1247 => x"66",
  1248 => x"66",
  1249 => x"66",
  1250 => x"3c",
  1251 => x"00",
  1252 => x"66",
  1253 => x"66",
  1254 => x"66",
  1255 => x"66",
  1256 => x"3c",
  1257 => x"3c",
  1258 => x"18",
  1259 => x"00",
  1260 => x"c6",
  1261 => x"c6",
  1262 => x"c6",
  1263 => x"d6",
  1264 => x"fe",
  1265 => x"ee",
  1266 => x"c6",
  1267 => x"00",
  1268 => x"c3",
  1269 => x"66",
  1270 => x"3c",
  1271 => x"18",
  1272 => x"3c",
  1273 => x"66",
  1274 => x"c3",
  1275 => x"00",
  1276 => x"c3",
  1277 => x"66",
  1278 => x"3c",
  1279 => x"18",
  1280 => x"18",
  1281 => x"18",
  1282 => x"18",
  1283 => x"00",
  1284 => x"fe",
  1285 => x"0c",
  1286 => x"18",
  1287 => x"30",
  1288 => x"60",
  1289 => x"c0",
  1290 => x"fe",
  1291 => x"00",
  1292 => x"3c",
  1293 => x"30",
  1294 => x"30",
  1295 => x"30",
  1296 => x"30",
  1297 => x"30",
  1298 => x"3c",
  1299 => x"00",
  1300 => x"c0",
  1301 => x"60",
  1302 => x"30",
  1303 => x"18",
  1304 => x"0c",
  1305 => x"06",
  1306 => x"03",
  1307 => x"00",
  1308 => x"3c",
  1309 => x"0c",
  1310 => x"0c",
  1311 => x"0c",
  1312 => x"0c",
  1313 => x"0c",
  1314 => x"3c",
  1315 => x"00",
  1316 => x"10",
  1317 => x"38",
  1318 => x"6c",
  1319 => x"c6",
  1320 => x"00",
  1321 => x"00",
  1322 => x"00",
  1323 => x"00",
  1324 => x"00",
  1325 => x"00",
  1326 => x"00",
  1327 => x"00",
  1328 => x"00",
  1329 => x"00",
  1330 => x"00",
  1331 => x"fe",
  1332 => x"18",
  1333 => x"18",
  1334 => x"0c",
  1335 => x"00",
  1336 => x"00",
  1337 => x"00",
  1338 => x"00",
  1339 => x"00",
  1340 => x"00",
  1341 => x"00",
  1342 => x"3c",
  1343 => x"06",
  1344 => x"3e",
  1345 => x"66",
  1346 => x"3e",
  1347 => x"00",
  1348 => x"60",
  1349 => x"60",
  1350 => x"7c",
  1351 => x"66",
  1352 => x"66",
  1353 => x"66",
  1354 => x"7c",
  1355 => x"00",
  1356 => x"00",
  1357 => x"00",
  1358 => x"3c",
  1359 => x"60",
  1360 => x"60",
  1361 => x"60",
  1362 => x"3c",
  1363 => x"00",
  1364 => x"06",
  1365 => x"06",
  1366 => x"3e",
  1367 => x"66",
  1368 => x"66",
  1369 => x"66",
  1370 => x"3e",
  1371 => x"00",
  1372 => x"00",
  1373 => x"00",
  1374 => x"3c",
  1375 => x"66",
  1376 => x"7e",
  1377 => x"60",
  1378 => x"3c",
  1379 => x"00",
  1380 => x"1c",
  1381 => x"30",
  1382 => x"7c",
  1383 => x"30",
  1384 => x"30",
  1385 => x"30",
  1386 => x"30",
  1387 => x"00",
  1388 => x"00",
  1389 => x"00",
  1390 => x"3e",
  1391 => x"66",
  1392 => x"66",
  1393 => x"3e",
  1394 => x"06",
  1395 => x"3c",
  1396 => x"60",
  1397 => x"60",
  1398 => x"7c",
  1399 => x"66",
  1400 => x"66",
  1401 => x"66",
  1402 => x"66",
  1403 => x"00",
  1404 => x"18",
  1405 => x"00",
  1406 => x"18",
  1407 => x"18",
  1408 => x"18",
  1409 => x"18",
  1410 => x"0c",
  1411 => x"00",
  1412 => x"0c",
  1413 => x"00",
  1414 => x"0c",
  1415 => x"0c",
  1416 => x"0c",
  1417 => x"0c",
  1418 => x"0c",
  1419 => x"78",
  1420 => x"60",
  1421 => x"60",
  1422 => x"66",
  1423 => x"6c",
  1424 => x"78",
  1425 => x"6c",
  1426 => x"66",
  1427 => x"00",
  1428 => x"18",
  1429 => x"18",
  1430 => x"18",
  1431 => x"18",
  1432 => x"18",
  1433 => x"18",
  1434 => x"0c",
  1435 => x"00",
  1436 => x"00",
  1437 => x"00",
  1438 => x"ec",
  1439 => x"fe",
  1440 => x"d6",
  1441 => x"c6",
  1442 => x"c6",
  1443 => x"00",
  1444 => x"00",
  1445 => x"00",
  1446 => x"7c",
  1447 => x"66",
  1448 => x"66",
  1449 => x"66",
  1450 => x"66",
  1451 => x"00",
  1452 => x"00",
  1453 => x"00",
  1454 => x"3c",
  1455 => x"66",
  1456 => x"66",
  1457 => x"66",
  1458 => x"3c",
  1459 => x"00",
  1460 => x"00",
  1461 => x"00",
  1462 => x"7c",
  1463 => x"66",
  1464 => x"66",
  1465 => x"7c",
  1466 => x"60",
  1467 => x"60",
  1468 => x"00",
  1469 => x"00",
  1470 => x"3e",
  1471 => x"66",
  1472 => x"66",
  1473 => x"3e",
  1474 => x"06",
  1475 => x"06",
  1476 => x"00",
  1477 => x"00",
  1478 => x"7c",
  1479 => x"66",
  1480 => x"60",
  1481 => x"60",
  1482 => x"60",
  1483 => x"00",
  1484 => x"00",
  1485 => x"00",
  1486 => x"3c",
  1487 => x"60",
  1488 => x"3c",
  1489 => x"06",
  1490 => x"7c",
  1491 => x"00",
  1492 => x"30",
  1493 => x"30",
  1494 => x"7c",
  1495 => x"30",
  1496 => x"30",
  1497 => x"30",
  1498 => x"1c",
  1499 => x"00",
  1500 => x"00",
  1501 => x"00",
  1502 => x"66",
  1503 => x"66",
  1504 => x"66",
  1505 => x"66",
  1506 => x"3e",
  1507 => x"00",
  1508 => x"00",
  1509 => x"00",
  1510 => x"66",
  1511 => x"66",
  1512 => x"66",
  1513 => x"3c",
  1514 => x"18",
  1515 => x"00",
  1516 => x"00",
  1517 => x"00",
  1518 => x"c6",
  1519 => x"c6",
  1520 => x"d6",
  1521 => x"fe",
  1522 => x"6c",
  1523 => x"00",
  1524 => x"00",
  1525 => x"00",
  1526 => x"c6",
  1527 => x"6c",
  1528 => x"38",
  1529 => x"6c",
  1530 => x"c6",
  1531 => x"00",
  1532 => x"00",
  1533 => x"00",
  1534 => x"66",
  1535 => x"66",
  1536 => x"66",
  1537 => x"3c",
  1538 => x"18",
  1539 => x"30",
  1540 => x"00",
  1541 => x"00",
  1542 => x"7e",
  1543 => x"0c",
  1544 => x"18",
  1545 => x"30",
  1546 => x"7e",
  1547 => x"00",
  1548 => x"0e",
  1549 => x"18",
  1550 => x"18",
  1551 => x"70",
  1552 => x"18",
  1553 => x"18",
  1554 => x"0e",
  1555 => x"00",
  1556 => x"18",
  1557 => x"18",
  1558 => x"18",
  1559 => x"18",
  1560 => x"18",
  1561 => x"18",
  1562 => x"18",
  1563 => x"00",
  1564 => x"70",
  1565 => x"18",
  1566 => x"18",
  1567 => x"0e",
  1568 => x"18",
  1569 => x"18",
  1570 => x"70",
  1571 => x"00",
  1572 => x"72",
  1573 => x"9c",
  1574 => x"00",
  1575 => x"00",
  1576 => x"00",
  1577 => x"00",
  1578 => x"00",
  1579 => x"00",
  1580 => x"fe",
  1581 => x"fe",
  1582 => x"fe",
  1583 => x"fe",
  1584 => x"fe",
  1585 => x"fe",
  1586 => x"fe",
  1587 => x"00",
  1588 => x"0a",
  1589 => x"0a",
  1590 => x"41",
  1591 => x"67",
  1592 => x"6e",
  1593 => x"75",
  1594 => x"73",
  1595 => x"20",
  1596 => x"49",
  1597 => x"44",
  1598 => x"3a",
  1599 => x"20",
  1600 => x"24",
  1601 => x"00",
  1602 => x"20",
  1603 => x"28",
  1604 => x"50",
  1605 => x"41",
  1606 => x"4c",
  1607 => x"29",
  1608 => x"00",
  1609 => x"20",
  1610 => x"28",
  1611 => x"4e",
  1612 => x"54",
  1613 => x"53",
  1614 => x"43",
  1615 => x"29",
  1616 => x"00",
  1617 => x"20",
  1618 => x"44",
  1619 => x"65",
  1620 => x"6e",
  1621 => x"69",
  1622 => x"73",
  1623 => x"65",
  1624 => x"20",
  1625 => x"49",
  1626 => x"44",
  1627 => x"3a",
  1628 => x"20",
  1629 => x"24",
  1630 => x"00",
  1631 => x"4d",
  1632 => x"65",
  1633 => x"6d",
  1634 => x"6f",
  1635 => x"72",
  1636 => x"79",
  1637 => x"20",
  1638 => x"62",
  1639 => x"61",
  1640 => x"73",
  1641 => x"65",
  1642 => x"3a",
  1643 => x"20",
  1644 => x"24",
  1645 => x"00",
  1646 => x"2c",
  1647 => x"20",
  1648 => x"73",
  1649 => x"69",
  1650 => x"7a",
  1651 => x"65",
  1652 => x"3a",
  1653 => x"20",
  1654 => x"24",
  1655 => x"00",
  1656 => x"5b",
  1657 => x"5f",
  1658 => x"5f",
  1659 => x"5f",
  1660 => x"5f",
  1661 => x"5f",
  1662 => x"5f",
  1663 => x"5f",
  1664 => x"5f",
  1665 => x"5f",
  1666 => x"5f",
  1667 => x"5f",
  1668 => x"5f",
  1669 => x"5f",
  1670 => x"5f",
  1671 => x"5f",
  1672 => x"5f",
  1673 => x"5f",
  1674 => x"5f",
  1675 => x"5f",
  1676 => x"5f",
  1677 => x"5f",
  1678 => x"5f",
  1679 => x"5f",
  1680 => x"5f",
  1681 => x"5f",
  1682 => x"5f",
  1683 => x"5f",
  1684 => x"5f",
  1685 => x"5f",
  1686 => x"5f",
  1687 => x"5f",
  1688 => x"5f",
  1689 => x"5d",
  1690 => x"00",
  1691 => x"0a",
  1692 => x"49",
  1693 => x"6e",
  1694 => x"63",
  1695 => x"6f",
  1696 => x"6d",
  1697 => x"70",
  1698 => x"61",
  1699 => x"74",
  1700 => x"69",
  1701 => x"62",
  1702 => x"6c",
  1703 => x"65",
  1704 => x"20",
  1705 => x"4d",
  1706 => x"65",
  1707 => x"6e",
  1708 => x"75",
  1709 => x"65",
  1710 => x"20",
  1711 => x"66",
  1712 => x"69",
  1713 => x"72",
  1714 => x"6d",
  1715 => x"77",
  1716 => x"61",
  1717 => x"72",
  1718 => x"65",
  1719 => x"21",
  1720 => x"00",
  1721 => x"0a",
  1722 => x"55",
  1723 => x"6e",
  1724 => x"6b",
  1725 => x"6e",
  1726 => x"6f",
  1727 => x"77",
  1728 => x"6e",
  1729 => x"20",
  1730 => x"63",
  1731 => x"6f",
  1732 => x"6d",
  1733 => x"6d",
  1734 => x"61",
  1735 => x"6e",
  1736 => x"64",
  1737 => x"3a",
  1738 => x"20",
  1739 => x"24",
  1740 => x"00",
  1741 => x"4d",
  1742 => x"69",
  1743 => x"6e",
  1744 => x"69",
  1745 => x"6d",
  1746 => x"69",
  1747 => x"67",
  1748 => x"20",
  1749 => x"62",
  1750 => x"79",
  1751 => x"20",
  1752 => x"44",
  1753 => x"65",
  1754 => x"6e",
  1755 => x"6e",
  1756 => x"69",
  1757 => x"73",
  1758 => x"20",
  1759 => x"76",
  1760 => x"61",
  1761 => x"6e",
  1762 => x"20",
  1763 => x"57",
  1764 => x"65",
  1765 => x"65",
  1766 => x"72",
  1767 => x"65",
  1768 => x"6e",
  1769 => x"20",
  1770 => x"0a",
  1771 => x"42",
  1772 => x"75",
  1773 => x"67",
  1774 => x"20",
  1775 => x"66",
  1776 => x"69",
  1777 => x"78",
  1778 => x"65",
  1779 => x"73",
  1780 => x"2c",
  1781 => x"20",
  1782 => x"6d",
  1783 => x"6f",
  1784 => x"64",
  1785 => x"73",
  1786 => x"20",
  1787 => x"61",
  1788 => x"6e",
  1789 => x"64",
  1790 => x"20",
  1791 => x"65",
  1792 => x"78",
  1793 => x"74",
  1794 => x"65",
  1795 => x"6e",
  1796 => x"73",
  1797 => x"69",
  1798 => x"6f",
  1799 => x"6e",
  1800 => x"73",
  1801 => x"20",
  1802 => x"62",
  1803 => x"79",
  1804 => x"20",
  1805 => x"4a",
  1806 => x"61",
  1807 => x"6b",
  1808 => x"75",
  1809 => x"62",
  1810 => x"20",
  1811 => x"42",
  1812 => x"65",
  1813 => x"64",
  1814 => x"6e",
  1815 => x"61",
  1816 => x"72",
  1817 => x"73",
  1818 => x"6b",
  1819 => x"69",
  1820 => x"20",
  1821 => x"61",
  1822 => x"6e",
  1823 => x"64",
  1824 => x"20",
  1825 => x"53",
  1826 => x"61",
  1827 => x"73",
  1828 => x"63",
  1829 => x"68",
  1830 => x"61",
  1831 => x"20",
  1832 => x"42",
  1833 => x"6f",
  1834 => x"69",
  1835 => x"6e",
  1836 => x"67",
  1837 => x"20",
  1838 => x"0a",
  1839 => x"54",
  1840 => x"47",
  1841 => x"36",
  1842 => x"38",
  1843 => x"4b",
  1844 => x"2e",
  1845 => x"43",
  1846 => x"20",
  1847 => x"28",
  1848 => x"36",
  1849 => x"38",
  1850 => x"30",
  1851 => x"30",
  1852 => x"30",
  1853 => x"20",
  1854 => x"49",
  1855 => x"50",
  1856 => x"20",
  1857 => x"43",
  1858 => x"6f",
  1859 => x"72",
  1860 => x"65",
  1861 => x"29",
  1862 => x"20",
  1863 => x"61",
  1864 => x"6e",
  1865 => x"64",
  1866 => x"20",
  1867 => x"43",
  1868 => x"68",
  1869 => x"61",
  1870 => x"6d",
  1871 => x"65",
  1872 => x"6c",
  1873 => x"65",
  1874 => x"6f",
  1875 => x"6e",
  1876 => x"20",
  1877 => x"50",
  1878 => x"6f",
  1879 => x"72",
  1880 => x"74",
  1881 => x"20",
  1882 => x"62",
  1883 => x"79",
  1884 => x"20",
  1885 => x"54",
  1886 => x"6f",
  1887 => x"62",
  1888 => x"69",
  1889 => x"61",
  1890 => x"73",
  1891 => x"20",
  1892 => x"47",
  1893 => x"75",
  1894 => x"62",
  1895 => x"65",
  1896 => x"6e",
  1897 => x"65",
  1898 => x"72",
  1899 => x"0a",
  1900 => x"00",
  1901 => x"0a",
  1902 => x"42",
  1903 => x"6f",
  1904 => x"6f",
  1905 => x"74",
  1906 => x"6c",
  1907 => x"6f",
  1908 => x"61",
  1909 => x"64",
  1910 => x"65",
  1911 => x"72",
  1912 => x"20",
  1913 => x"20",
  1914 => x"20",
  1915 => x"20",
  1916 => x"32",
  1917 => x"30",
  1918 => x"31",
  1919 => x"30",
  1920 => x"2d",
  1921 => x"30",
  1922 => x"39",
  1923 => x"2d",
  1924 => x"31",
  1925 => x"30",
  1926 => x"00",
  1927 => x"0a",
  1928 => x"4d",
  1929 => x"69",
  1930 => x"6e",
  1931 => x"69",
  1932 => x"6d",
  1933 => x"69",
  1934 => x"67",
  1935 => x"20",
  1936 => x"63",
  1937 => x"6f",
  1938 => x"72",
  1939 => x"65",
  1940 => x"20",
  1941 => x"20",
  1942 => x"32",
  1943 => x"30",
  1944 => x"31",
  1945 => x"31",
  1946 => x"2d",
  1947 => x"30",
  1948 => x"34",
  1949 => x"2d",
  1950 => x"31",
  1951 => x"30",
  1952 => x"00",
	others => x"00"
);

begin

-- We use a dual-port RAM here - one port for the lower byte, one for the upper byte.  This allows us to
-- present a 16-bit interface while allowing byte writes.

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and lds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1'))) := d(7 downto 0);
			q(7 downto 0) <= d(7 downto 0);
		else
			q(7 downto 0) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'1')));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if we_n = '0' and uds_n='0' then
			ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0'))) := d(15 downto 8);
			q(15 downto 8) <= d(15 downto 8);
		else
			q(15 downto 8) <= ram(to_integer(unsigned(addr(maxAddrBitBRAM downto 1)&'0')));
		end if;
	end if;
end process;

end arch;

